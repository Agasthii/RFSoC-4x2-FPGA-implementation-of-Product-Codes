`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/11/2024 07:25:58 AM
// Design Name: 
// Module Name: PC_datapath_ebch_256_239_new
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PC_datapath_testing #(
    parameter k = 239,
    parameter n = 256,
    parameter depth = 16
    )(
    input wire clk,
    input wire reset,
    input wire [4095:0] seed,
    input wire [15:0] cross_prob,
    input wire [4:0] iterations,
    output reg [63:0] errs,
    output reg [63:0] errs_u,
//    output reg [63:0] errs_u,
    output reg [63:0] sims
    );
    
    wire new;
    wire hold_enc;
    wire store; // store out_codewords from the encoder
    
    reg uncoded; // for uncoded error calculation
    reg [3:0] uncoded_last_iter; // the last set of the uncoded error calculation. Here we only consider 15 not 16
    
    wire [n-1:0] codeword1;
    wire [n-1:0] codeword2;
    wire [n-1:0] codeword3;
    wire [n-1:0] codeword4;
    wire [n-1:0] codeword5;
    wire [n-1:0] codeword6;
    wire [n-1:0] codeword7;
    wire [n-1:0] codeword8;
    wire [n-1:0] codeword9;
    wire [n-1:0] codeword10;
    wire [n-1:0] codeword11;
    wire [n-1:0] codeword12;
    wire [n-1:0] codeword13;
    wire [n-1:0] codeword14;
    wire [n-1:0] codeword15;
    wire [n-1:0] codeword16; 
    
    PC_encoding_block_testing PC_encoding_block_testing_d(
        .clk(clk),
        .reset(reset),
        .seed(seed),
        .new1(new),
        .hold_enc(hold_enc),
        .store(store),
        .out_codeword1(codeword1),
        .out_codeword2(codeword2),
        .out_codeword3(codeword3),
        .out_codeword4(codeword4),
        .out_codeword5(codeword5),
        .out_codeword6(codeword6),
        .out_codeword7(codeword7),
        .out_codeword8(codeword8),
        .out_codeword9(codeword9),
        .out_codeword10(codeword10),
        .out_codeword11(codeword11),
        .out_codeword12(codeword12),
        .out_codeword13(codeword13),
        .out_codeword14(codeword14),
        .out_codeword15(codeword15),
        .out_codeword16(codeword16)
        );
        
    wire [n-1:0] received1;
    wire [n-1:0] received2;
    wire [n-1:0] received3;
    wire [n-1:0] received4;
    wire [n-1:0] received5;
    wire [n-1:0] received6;
    wire [n-1:0] received7;
    wire [n-1:0] received8;
    wire [n-1:0] received9;
    wire [n-1:0] received10;
    wire [n-1:0] received11;
    wire [n-1:0] received12;
    wire [n-1:0] received13;
    wire [n-1:0] received14;
    wire [n-1:0] received15;
    wire [n-1:0] received16;
        
    PC_bsc_channel_block_ebch_256_239 PC_bsc_channel_block_ebch_256_239_d(
        .clk(clk),
        .reset(reset),
        .seed(seed),
        .cross_prob(cross_prob),
        .codeword1(codeword1),
        .codeword2(codeword2),
        .codeword3(codeword3),
        .codeword4(codeword4),
        .codeword5(codeword5),
        .codeword6(codeword6),
        .codeword7(codeword7),
        .codeword8(codeword8),
        .codeword9(codeword9),
        .codeword10(codeword10),
        .codeword11(codeword11),
        .codeword12(codeword12),
        .codeword13(codeword13),
        .codeword14(codeword14),
        .codeword15(codeword15),
        .codeword16(codeword16),
        .received1(received1),
        .received2(received2),
        .received3(received3),
        .received4(received4),
        .received5(received5),
        .received6(received6),
        .received7(received7),
        .received8(received8),
        .received9(received9),
        .received10(received10),
        .received11(received11),
        .received12(received12),
        .received13(received13),
        .received14(received14),
        .received15(received15),
        .received16(received16)
        );
        
    wire valid1;
    wire valid2;
    wire valid_err;
    
    wire [n-1:0] dec1;
    wire [n-1:0] dec2;
    wire [n-1:0] dec3;
    wire [n-1:0] dec4;
    wire [n-1:0] dec5;
    wire [n-1:0] dec6;
    wire [n-1:0] dec7;
    wire [n-1:0] dec8;
    wire [n-1:0] dec9;
    wire [n-1:0] dec10;
    wire [n-1:0] dec11;
    wire [n-1:0] dec12;
    wire [n-1:0] dec13;
    wire [n-1:0] dec14;
    wire [n-1:0] dec15;
    wire [n-1:0] dec16;
        
    PC_decoding_block_ebch_256_239 PC_decoding_block_ebch_256_239_d(
        .clk(clk),
        .reset(reset),
        .new(new),
        .hold_enc(hold_enc),
        .iter(iterations),
        .rec1(received1),
        .rec2(received2),
        .rec3(received3),
        .rec4(received4),
        .rec5(received5),
        .rec6(received6),
        .rec7(received7),
        .rec8(received8),
        .rec9(received9),
        .rec10(received10),
        .rec11(received11),
        .rec12(received12),
        .rec13(received13),
        .rec14(received14),
        .rec15(received15),
        .rec16(received16),
        .valid1(valid1),
        .valid2(valid2),
        .valid_err(valid_err),
        .dec1(dec1),
        .dec2(dec2),
        .dec3(dec3),
        .dec4(dec4),
        .dec5(dec5),
        .dec6(dec6),
        .dec7(dec7),
        .dec8(dec8),
        .dec9(dec9),
        .dec10(dec10),
        .dec11(dec11),
        .dec12(dec12),
        .dec13(dec13),
        .dec14(dec14),
        .dec15(dec15),
        .dec16(dec16)
        );
        
    reg [9:0] fifo_depth;
    
    reg [4:0] x;
    
    reg valid_err_count = 1'b0;
    reg valid_err_sum = 1'b0;
    
    // For the encoded codewords
    reg [(16*n-1):0] FIFO_1;
    reg [(16*n-1):0] FIFO_2;
    reg [(16*n-1):0] FIFO_3;
    reg [(16*n-1):0] FIFO_4;
    reg [(16*n-1):0] FIFO_5;
    reg [(16*n-1):0] FIFO_6;
    reg [(16*n-1):0] FIFO_7;
    reg [(16*n-1):0] FIFO_8;
    reg [(16*n-1):0] FIFO_9;
    reg [(16*n-1):0] FIFO_10;
    reg [(16*n-1):0] FIFO_11;
    reg [(16*n-1):0] FIFO_12;
    reg [(16*n-1):0] FIFO_13;
    reg [(16*n-1):0] FIFO_14;
    reg [(16*n-1):0] FIFO_15;
    reg [(16*n-1):0] FIFO_16;
    
    reg [(n-1):0] error_vector1;
    reg [(n-1):0] error_vector2;
    reg [(n-1):0] error_vector3;
    reg [(n-1):0] error_vector4;
    reg [(n-1):0] error_vector5;
    reg [(n-1):0] error_vector6;
    reg [(n-1):0] error_vector7;
    reg [(n-1):0] error_vector8;
    reg [(n-1):0] error_vector9;
    reg [(n-1):0] error_vector10;
    reg [(n-1):0] error_vector11;
    reg [(n-1):0] error_vector12;
    reg [(n-1):0] error_vector13;
    reg [(n-1):0] error_vector14;
    reg [(n-1):0] error_vector15;
    reg [(n-1):0] error_vector16;
    
    reg [8:0] errs1;
    reg [8:0] errs2;
    reg [8:0] errs3;
    reg [8:0] errs4;
    reg [8:0] errs5;
    reg [8:0] errs6;
    reg [8:0] errs7;
    reg [8:0] errs8;
    reg [8:0] errs9;
    reg [8:0] errs10;
    reg [8:0] errs11;
    reg [8:0] errs12;
    reg [8:0] errs13;
    reg [8:0] errs14;
    reg [8:0] errs15;
    reg [8:0] errs16;


    // Uncoded errors
    reg [(n-1):0] error_u_vector1;
    reg [(n-1):0] error_u_vector2;
    reg [(n-1):0] error_u_vector3;
    reg [(n-1):0] error_u_vector4;
    reg [(n-1):0] error_u_vector5;
    reg [(n-1):0] error_u_vector6;
    reg [(n-1):0] error_u_vector7;
    reg [(n-1):0] error_u_vector8;
    reg [(n-1):0] error_u_vector9;
    reg [(n-1):0] error_u_vector10;
    reg [(n-1):0] error_u_vector11;
    reg [(n-1):0] error_u_vector12;
    reg [(n-1):0] error_u_vector13;
    reg [(n-1):0] error_u_vector14;
    reg [(n-1):0] error_u_vector15;
    reg [(n-1):0] error_u_vector16;
    
    reg [8:0] errs1_u;
    reg [8:0] errs2_u;
    reg [8:0] errs3_u;
    reg [8:0] errs4_u;
    reg [8:0] errs5_u;
    reg [8:0] errs6_u;
    reg [8:0] errs7_u;
    reg [8:0] errs8_u;
    reg [8:0] errs9_u;
    reg [8:0] errs10_u;
    reg [8:0] errs11_u;
    reg [8:0] errs12_u;
    reg [8:0] errs13_u;
    reg [8:0] errs14_u;
    reg [8:0] errs15_u;
    reg [8:0] errs16_u;
    
    reg counting;
    
    integer i;
    
    always@(posedge clk) begin
        if(reset) begin
        
            if (store) begin

                uncoded <= 1'b1;
                uncoded_last_iter <= uncoded_last_iter + 4'b1;
                
                // Shift the FIFO buffer
                FIFO_1 <= (FIFO_1 << n);
                FIFO_2 <= (FIFO_2 << n);
                FIFO_3 <= (FIFO_3 << n);
                FIFO_4 <= (FIFO_4 << n);
                FIFO_5 <= (FIFO_5 << n);
                FIFO_6 <= (FIFO_6 << n);
                FIFO_7 <= (FIFO_7 << n);
                FIFO_8 <= (FIFO_8 << n);
                FIFO_9 <= (FIFO_9 << n);
                FIFO_10 <= (FIFO_10 << n);
                FIFO_11 <= (FIFO_11 << n);
                FIFO_12 <= (FIFO_12 << n);
                FIFO_13 <= (FIFO_13 << n);
                FIFO_14 <= (FIFO_14 << n);
                FIFO_15 <= (FIFO_15 << n);
                FIFO_16 <= (FIFO_16 << n);
                
                // Store the new codeword in the FIFO
                FIFO_1[(n-1):0] <= codeword1;
                FIFO_2[(n-1):0] <= codeword2;
                FIFO_3[(n-1):0] <= codeword3;
                FIFO_4[(n-1):0] <= codeword4;
                FIFO_5[(n-1):0] <= codeword5;
                FIFO_6[(n-1):0] <= codeword6;
                FIFO_7[(n-1):0] <= codeword7;
                FIFO_8[(n-1):0] <= codeword8;
                FIFO_9[(n-1):0] <= codeword9;
                FIFO_10[(n-1):0] <= codeword10;
                FIFO_11[(n-1):0] <= codeword11;
                FIFO_12[(n-1):0] <= codeword12;
                FIFO_13[(n-1):0] <= codeword13;
                FIFO_14[(n-1):0] <= codeword14;
                FIFO_15[(n-1):0] <= codeword15;
                FIFO_16[(n-1):0] <= codeword16;

            end else begin
                uncoded <= 1'b0;
                uncoded_last_iter <= 4'b0;
            end

            if ((uncoded)&(store)) begin
                //Uncoded error vectors
                error_u_vector1 <= FIFO_1[(n-1):0] ^ received1; 
                error_u_vector2 <= FIFO_2[(n-1):0] ^ received2; 
                error_u_vector3 <= FIFO_3[(n-1):0] ^ received3; 
                error_u_vector4 <= FIFO_4[(n-1):0] ^ received4; 
                error_u_vector5 <= FIFO_5[(n-1):0] ^ received5; 
                error_u_vector6 <= FIFO_6[(n-1):0] ^ received6; 
                error_u_vector7 <= FIFO_7[(n-1):0] ^ received7; 
                error_u_vector8 <= FIFO_8[(n-1):0] ^ received8; 
                error_u_vector9 <= FIFO_9[(n-1):0] ^ received9; 
                error_u_vector10 <= FIFO_10[(n-1):0] ^ received10; 
                error_u_vector11 <= FIFO_11[(n-1):0] ^ received11; 
                error_u_vector12 <= FIFO_12[(n-1):0] ^ received12; 
                error_u_vector13 <= FIFO_13[(n-1):0] ^ received13; 
                error_u_vector14 <= FIFO_14[(n-1):0] ^ received14; 
                error_u_vector15 <= FIFO_15[(n-1):0] ^ received15; 
                error_u_vector16 <= FIFO_16[(n-1):0] ^ received16; 

            end else begin
                error_u_vector1 <= 0;
                error_u_vector2 <= 0;
                error_u_vector3 <= 0;
                error_u_vector4 <= 0;
                error_u_vector5 <= 0;
                error_u_vector6 <= 0;
                error_u_vector7 <= 0;
                error_u_vector8 <= 0;
                error_u_vector9 <= 0;
                error_u_vector10 <= 0;
                error_u_vector11 <= 0;
                error_u_vector12 <= 0;
                error_u_vector13 <= 0;
                error_u_vector14 <= 0;
                error_u_vector15 <= 0;
                error_u_vector16 <= 0;

            end
            
            if (valid2) begin
                x <= x + 1;
            
                error_vector1 <= dec1 ^ {FIFO_16[256*0+x*16+0],FIFO_15[256*0+x*16+0],FIFO_14[256*0+x*16+0],FIFO_13[256*0+x*16+0],FIFO_12[256*0+x*16+0],FIFO_11[256*0+x*16+0],FIFO_10[256*0+x*16+0],FIFO_9[256*0+x*16+0],FIFO_8[256*0+x*16+0],FIFO_7[256*0+x*16+0],FIFO_6[256*0+x*16+0],FIFO_5[256*0+x*16+0],FIFO_4[256*0+x*16+0],FIFO_3[256*0+x*16+0],FIFO_2[256*0+x*16+0],FIFO_1[256*0+x*16+0],FIFO_16[256*1+x*16+0],FIFO_15[256*1+x*16+0],FIFO_14[256*1+x*16+0],FIFO_13[256*1+x*16+0],FIFO_12[256*1+x*16+0],FIFO_11[256*1+x*16+0],FIFO_10[256*1+x*16+0],FIFO_9[256*1+x*16+0],FIFO_8[256*1+x*16+0],FIFO_7[256*1+x*16+0],FIFO_6[256*1+x*16+0],FIFO_5[256*1+x*16+0],FIFO_4[256*1+x*16+0],FIFO_3[256*1+x*16+0],FIFO_2[256*1+x*16+0],FIFO_1[256*1+x*16+0],FIFO_16[256*2+x*16+0],FIFO_15[256*2+x*16+0],FIFO_14[256*2+x*16+0],FIFO_13[256*2+x*16+0],FIFO_12[256*2+x*16+0],FIFO_11[256*2+x*16+0],FIFO_10[256*2+x*16+0],FIFO_9[256*2+x*16+0],FIFO_8[256*2+x*16+0],FIFO_7[256*2+x*16+0],FIFO_6[256*2+x*16+0],FIFO_5[256*2+x*16+0],FIFO_4[256*2+x*16+0],FIFO_3[256*2+x*16+0],FIFO_2[256*2+x*16+0],FIFO_1[256*2+x*16+0],FIFO_16[256*3+x*16+0],FIFO_15[256*3+x*16+0],FIFO_14[256*3+x*16+0],FIFO_13[256*3+x*16+0],FIFO_12[256*3+x*16+0],FIFO_11[256*3+x*16+0],FIFO_10[256*3+x*16+0],FIFO_9[256*3+x*16+0],FIFO_8[256*3+x*16+0],FIFO_7[256*3+x*16+0],FIFO_6[256*3+x*16+0],FIFO_5[256*3+x*16+0],FIFO_4[256*3+x*16+0],FIFO_3[256*3+x*16+0],FIFO_2[256*3+x*16+0],FIFO_1[256*3+x*16+0],FIFO_16[256*4+x*16+0],FIFO_15[256*4+x*16+0],FIFO_14[256*4+x*16+0],FIFO_13[256*4+x*16+0],FIFO_12[256*4+x*16+0],FIFO_11[256*4+x*16+0],FIFO_10[256*4+x*16+0],FIFO_9[256*4+x*16+0],FIFO_8[256*4+x*16+0],FIFO_7[256*4+x*16+0],FIFO_6[256*4+x*16+0],FIFO_5[256*4+x*16+0],FIFO_4[256*4+x*16+0],FIFO_3[256*4+x*16+0],FIFO_2[256*4+x*16+0],FIFO_1[256*4+x*16+0],FIFO_16[256*5+x*16+0],FIFO_15[256*5+x*16+0],FIFO_14[256*5+x*16+0],FIFO_13[256*5+x*16+0],FIFO_12[256*5+x*16+0],FIFO_11[256*5+x*16+0],FIFO_10[256*5+x*16+0],FIFO_9[256*5+x*16+0],FIFO_8[256*5+x*16+0],FIFO_7[256*5+x*16+0],FIFO_6[256*5+x*16+0],FIFO_5[256*5+x*16+0],FIFO_4[256*5+x*16+0],FIFO_3[256*5+x*16+0],FIFO_2[256*5+x*16+0],FIFO_1[256*5+x*16+0],FIFO_16[256*6+x*16+0],FIFO_15[256*6+x*16+0],FIFO_14[256*6+x*16+0],FIFO_13[256*6+x*16+0],FIFO_12[256*6+x*16+0],FIFO_11[256*6+x*16+0],FIFO_10[256*6+x*16+0],FIFO_9[256*6+x*16+0],FIFO_8[256*6+x*16+0],FIFO_7[256*6+x*16+0],FIFO_6[256*6+x*16+0],FIFO_5[256*6+x*16+0],FIFO_4[256*6+x*16+0],FIFO_3[256*6+x*16+0],FIFO_2[256*6+x*16+0],FIFO_1[256*6+x*16+0],FIFO_16[256*7+x*16+0],FIFO_15[256*7+x*16+0],FIFO_14[256*7+x*16+0],FIFO_13[256*7+x*16+0],FIFO_12[256*7+x*16+0],FIFO_11[256*7+x*16+0],FIFO_10[256*7+x*16+0],FIFO_9[256*7+x*16+0],FIFO_8[256*7+x*16+0],FIFO_7[256*7+x*16+0],FIFO_6[256*7+x*16+0],FIFO_5[256*7+x*16+0],FIFO_4[256*7+x*16+0],FIFO_3[256*7+x*16+0],FIFO_2[256*7+x*16+0],FIFO_1[256*7+x*16+0],FIFO_16[256*8+x*16+0],FIFO_15[256*8+x*16+0],FIFO_14[256*8+x*16+0],FIFO_13[256*8+x*16+0],FIFO_12[256*8+x*16+0],FIFO_11[256*8+x*16+0],FIFO_10[256*8+x*16+0],FIFO_9[256*8+x*16+0],FIFO_8[256*8+x*16+0],FIFO_7[256*8+x*16+0],FIFO_6[256*8+x*16+0],FIFO_5[256*8+x*16+0],FIFO_4[256*8+x*16+0],FIFO_3[256*8+x*16+0],FIFO_2[256*8+x*16+0],FIFO_1[256*8+x*16+0],FIFO_16[256*9+x*16+0],FIFO_15[256*9+x*16+0],FIFO_14[256*9+x*16+0],FIFO_13[256*9+x*16+0],FIFO_12[256*9+x*16+0],FIFO_11[256*9+x*16+0],FIFO_10[256*9+x*16+0],FIFO_9[256*9+x*16+0],FIFO_8[256*9+x*16+0],FIFO_7[256*9+x*16+0],FIFO_6[256*9+x*16+0],FIFO_5[256*9+x*16+0],FIFO_4[256*9+x*16+0],FIFO_3[256*9+x*16+0],FIFO_2[256*9+x*16+0],FIFO_1[256*9+x*16+0],FIFO_16[256*10+x*16+0],FIFO_15[256*10+x*16+0],FIFO_14[256*10+x*16+0],FIFO_13[256*10+x*16+0],FIFO_12[256*10+x*16+0],FIFO_11[256*10+x*16+0],FIFO_10[256*10+x*16+0],FIFO_9[256*10+x*16+0],FIFO_8[256*10+x*16+0],FIFO_7[256*10+x*16+0],FIFO_6[256*10+x*16+0],FIFO_5[256*10+x*16+0],FIFO_4[256*10+x*16+0],FIFO_3[256*10+x*16+0],FIFO_2[256*10+x*16+0],FIFO_1[256*10+x*16+0],FIFO_16[256*11+x*16+0],FIFO_15[256*11+x*16+0],FIFO_14[256*11+x*16+0],FIFO_13[256*11+x*16+0],FIFO_12[256*11+x*16+0],FIFO_11[256*11+x*16+0],FIFO_10[256*11+x*16+0],FIFO_9[256*11+x*16+0],FIFO_8[256*11+x*16+0],FIFO_7[256*11+x*16+0],FIFO_6[256*11+x*16+0],FIFO_5[256*11+x*16+0],FIFO_4[256*11+x*16+0],FIFO_3[256*11+x*16+0],FIFO_2[256*11+x*16+0],FIFO_1[256*11+x*16+0],FIFO_16[256*12+x*16+0],FIFO_15[256*12+x*16+0],FIFO_14[256*12+x*16+0],FIFO_13[256*12+x*16+0],FIFO_12[256*12+x*16+0],FIFO_11[256*12+x*16+0],FIFO_10[256*12+x*16+0],FIFO_9[256*12+x*16+0],FIFO_8[256*12+x*16+0],FIFO_7[256*12+x*16+0],FIFO_6[256*12+x*16+0],FIFO_5[256*12+x*16+0],FIFO_4[256*12+x*16+0],FIFO_3[256*12+x*16+0],FIFO_2[256*12+x*16+0],FIFO_1[256*12+x*16+0],FIFO_16[256*13+x*16+0],FIFO_15[256*13+x*16+0],FIFO_14[256*13+x*16+0],FIFO_13[256*13+x*16+0],FIFO_12[256*13+x*16+0],FIFO_11[256*13+x*16+0],FIFO_10[256*13+x*16+0],FIFO_9[256*13+x*16+0],FIFO_8[256*13+x*16+0],FIFO_7[256*13+x*16+0],FIFO_6[256*13+x*16+0],FIFO_5[256*13+x*16+0],FIFO_4[256*13+x*16+0],FIFO_3[256*13+x*16+0],FIFO_2[256*13+x*16+0],FIFO_1[256*13+x*16+0],FIFO_16[256*14+x*16+0],FIFO_15[256*14+x*16+0],FIFO_14[256*14+x*16+0],FIFO_13[256*14+x*16+0],FIFO_12[256*14+x*16+0],FIFO_11[256*14+x*16+0],FIFO_10[256*14+x*16+0],FIFO_9[256*14+x*16+0],FIFO_8[256*14+x*16+0],FIFO_7[256*14+x*16+0],FIFO_6[256*14+x*16+0],FIFO_5[256*14+x*16+0],FIFO_4[256*14+x*16+0],FIFO_3[256*14+x*16+0],FIFO_2[256*14+x*16+0],FIFO_1[256*14+x*16+0],FIFO_16[256*15+x*16+0],FIFO_15[256*15+x*16+0],FIFO_14[256*15+x*16+0],FIFO_13[256*15+x*16+0],FIFO_12[256*15+x*16+0],FIFO_11[256*15+x*16+0],FIFO_10[256*15+x*16+0],FIFO_9[256*15+x*16+0],FIFO_8[256*15+x*16+0],FIFO_7[256*15+x*16+0],FIFO_6[256*15+x*16+0],FIFO_5[256*15+x*16+0],FIFO_4[256*15+x*16+0],FIFO_3[256*15+x*16+0],FIFO_2[256*15+x*16+0],FIFO_1[256*15+x*16+0]}; 
                error_vector2 <= dec2 ^ {FIFO_16[256*0+x*16+1],FIFO_15[256*0+x*16+1],FIFO_14[256*0+x*16+1],FIFO_13[256*0+x*16+1],FIFO_12[256*0+x*16+1],FIFO_11[256*0+x*16+1],FIFO_10[256*0+x*16+1],FIFO_9[256*0+x*16+1],FIFO_8[256*0+x*16+1],FIFO_7[256*0+x*16+1],FIFO_6[256*0+x*16+1],FIFO_5[256*0+x*16+1],FIFO_4[256*0+x*16+1],FIFO_3[256*0+x*16+1],FIFO_2[256*0+x*16+1],FIFO_1[256*0+x*16+1],FIFO_16[256*1+x*16+1],FIFO_15[256*1+x*16+1],FIFO_14[256*1+x*16+1],FIFO_13[256*1+x*16+1],FIFO_12[256*1+x*16+1],FIFO_11[256*1+x*16+1],FIFO_10[256*1+x*16+1],FIFO_9[256*1+x*16+1],FIFO_8[256*1+x*16+1],FIFO_7[256*1+x*16+1],FIFO_6[256*1+x*16+1],FIFO_5[256*1+x*16+1],FIFO_4[256*1+x*16+1],FIFO_3[256*1+x*16+1],FIFO_2[256*1+x*16+1],FIFO_1[256*1+x*16+1],FIFO_16[256*2+x*16+1],FIFO_15[256*2+x*16+1],FIFO_14[256*2+x*16+1],FIFO_13[256*2+x*16+1],FIFO_12[256*2+x*16+1],FIFO_11[256*2+x*16+1],FIFO_10[256*2+x*16+1],FIFO_9[256*2+x*16+1],FIFO_8[256*2+x*16+1],FIFO_7[256*2+x*16+1],FIFO_6[256*2+x*16+1],FIFO_5[256*2+x*16+1],FIFO_4[256*2+x*16+1],FIFO_3[256*2+x*16+1],FIFO_2[256*2+x*16+1],FIFO_1[256*2+x*16+1],FIFO_16[256*3+x*16+1],FIFO_15[256*3+x*16+1],FIFO_14[256*3+x*16+1],FIFO_13[256*3+x*16+1],FIFO_12[256*3+x*16+1],FIFO_11[256*3+x*16+1],FIFO_10[256*3+x*16+1],FIFO_9[256*3+x*16+1],FIFO_8[256*3+x*16+1],FIFO_7[256*3+x*16+1],FIFO_6[256*3+x*16+1],FIFO_5[256*3+x*16+1],FIFO_4[256*3+x*16+1],FIFO_3[256*3+x*16+1],FIFO_2[256*3+x*16+1],FIFO_1[256*3+x*16+1],FIFO_16[256*4+x*16+1],FIFO_15[256*4+x*16+1],FIFO_14[256*4+x*16+1],FIFO_13[256*4+x*16+1],FIFO_12[256*4+x*16+1],FIFO_11[256*4+x*16+1],FIFO_10[256*4+x*16+1],FIFO_9[256*4+x*16+1],FIFO_8[256*4+x*16+1],FIFO_7[256*4+x*16+1],FIFO_6[256*4+x*16+1],FIFO_5[256*4+x*16+1],FIFO_4[256*4+x*16+1],FIFO_3[256*4+x*16+1],FIFO_2[256*4+x*16+1],FIFO_1[256*4+x*16+1],FIFO_16[256*5+x*16+1],FIFO_15[256*5+x*16+1],FIFO_14[256*5+x*16+1],FIFO_13[256*5+x*16+1],FIFO_12[256*5+x*16+1],FIFO_11[256*5+x*16+1],FIFO_10[256*5+x*16+1],FIFO_9[256*5+x*16+1],FIFO_8[256*5+x*16+1],FIFO_7[256*5+x*16+1],FIFO_6[256*5+x*16+1],FIFO_5[256*5+x*16+1],FIFO_4[256*5+x*16+1],FIFO_3[256*5+x*16+1],FIFO_2[256*5+x*16+1],FIFO_1[256*5+x*16+1],FIFO_16[256*6+x*16+1],FIFO_15[256*6+x*16+1],FIFO_14[256*6+x*16+1],FIFO_13[256*6+x*16+1],FIFO_12[256*6+x*16+1],FIFO_11[256*6+x*16+1],FIFO_10[256*6+x*16+1],FIFO_9[256*6+x*16+1],FIFO_8[256*6+x*16+1],FIFO_7[256*6+x*16+1],FIFO_6[256*6+x*16+1],FIFO_5[256*6+x*16+1],FIFO_4[256*6+x*16+1],FIFO_3[256*6+x*16+1],FIFO_2[256*6+x*16+1],FIFO_1[256*6+x*16+1],FIFO_16[256*7+x*16+1],FIFO_15[256*7+x*16+1],FIFO_14[256*7+x*16+1],FIFO_13[256*7+x*16+1],FIFO_12[256*7+x*16+1],FIFO_11[256*7+x*16+1],FIFO_10[256*7+x*16+1],FIFO_9[256*7+x*16+1],FIFO_8[256*7+x*16+1],FIFO_7[256*7+x*16+1],FIFO_6[256*7+x*16+1],FIFO_5[256*7+x*16+1],FIFO_4[256*7+x*16+1],FIFO_3[256*7+x*16+1],FIFO_2[256*7+x*16+1],FIFO_1[256*7+x*16+1],FIFO_16[256*8+x*16+1],FIFO_15[256*8+x*16+1],FIFO_14[256*8+x*16+1],FIFO_13[256*8+x*16+1],FIFO_12[256*8+x*16+1],FIFO_11[256*8+x*16+1],FIFO_10[256*8+x*16+1],FIFO_9[256*8+x*16+1],FIFO_8[256*8+x*16+1],FIFO_7[256*8+x*16+1],FIFO_6[256*8+x*16+1],FIFO_5[256*8+x*16+1],FIFO_4[256*8+x*16+1],FIFO_3[256*8+x*16+1],FIFO_2[256*8+x*16+1],FIFO_1[256*8+x*16+1],FIFO_16[256*9+x*16+1],FIFO_15[256*9+x*16+1],FIFO_14[256*9+x*16+1],FIFO_13[256*9+x*16+1],FIFO_12[256*9+x*16+1],FIFO_11[256*9+x*16+1],FIFO_10[256*9+x*16+1],FIFO_9[256*9+x*16+1],FIFO_8[256*9+x*16+1],FIFO_7[256*9+x*16+1],FIFO_6[256*9+x*16+1],FIFO_5[256*9+x*16+1],FIFO_4[256*9+x*16+1],FIFO_3[256*9+x*16+1],FIFO_2[256*9+x*16+1],FIFO_1[256*9+x*16+1],FIFO_16[256*10+x*16+1],FIFO_15[256*10+x*16+1],FIFO_14[256*10+x*16+1],FIFO_13[256*10+x*16+1],FIFO_12[256*10+x*16+1],FIFO_11[256*10+x*16+1],FIFO_10[256*10+x*16+1],FIFO_9[256*10+x*16+1],FIFO_8[256*10+x*16+1],FIFO_7[256*10+x*16+1],FIFO_6[256*10+x*16+1],FIFO_5[256*10+x*16+1],FIFO_4[256*10+x*16+1],FIFO_3[256*10+x*16+1],FIFO_2[256*10+x*16+1],FIFO_1[256*10+x*16+1],FIFO_16[256*11+x*16+1],FIFO_15[256*11+x*16+1],FIFO_14[256*11+x*16+1],FIFO_13[256*11+x*16+1],FIFO_12[256*11+x*16+1],FIFO_11[256*11+x*16+1],FIFO_10[256*11+x*16+1],FIFO_9[256*11+x*16+1],FIFO_8[256*11+x*16+1],FIFO_7[256*11+x*16+1],FIFO_6[256*11+x*16+1],FIFO_5[256*11+x*16+1],FIFO_4[256*11+x*16+1],FIFO_3[256*11+x*16+1],FIFO_2[256*11+x*16+1],FIFO_1[256*11+x*16+1],FIFO_16[256*12+x*16+1],FIFO_15[256*12+x*16+1],FIFO_14[256*12+x*16+1],FIFO_13[256*12+x*16+1],FIFO_12[256*12+x*16+1],FIFO_11[256*12+x*16+1],FIFO_10[256*12+x*16+1],FIFO_9[256*12+x*16+1],FIFO_8[256*12+x*16+1],FIFO_7[256*12+x*16+1],FIFO_6[256*12+x*16+1],FIFO_5[256*12+x*16+1],FIFO_4[256*12+x*16+1],FIFO_3[256*12+x*16+1],FIFO_2[256*12+x*16+1],FIFO_1[256*12+x*16+1],FIFO_16[256*13+x*16+1],FIFO_15[256*13+x*16+1],FIFO_14[256*13+x*16+1],FIFO_13[256*13+x*16+1],FIFO_12[256*13+x*16+1],FIFO_11[256*13+x*16+1],FIFO_10[256*13+x*16+1],FIFO_9[256*13+x*16+1],FIFO_8[256*13+x*16+1],FIFO_7[256*13+x*16+1],FIFO_6[256*13+x*16+1],FIFO_5[256*13+x*16+1],FIFO_4[256*13+x*16+1],FIFO_3[256*13+x*16+1],FIFO_2[256*13+x*16+1],FIFO_1[256*13+x*16+1],FIFO_16[256*14+x*16+1],FIFO_15[256*14+x*16+1],FIFO_14[256*14+x*16+1],FIFO_13[256*14+x*16+1],FIFO_12[256*14+x*16+1],FIFO_11[256*14+x*16+1],FIFO_10[256*14+x*16+1],FIFO_9[256*14+x*16+1],FIFO_8[256*14+x*16+1],FIFO_7[256*14+x*16+1],FIFO_6[256*14+x*16+1],FIFO_5[256*14+x*16+1],FIFO_4[256*14+x*16+1],FIFO_3[256*14+x*16+1],FIFO_2[256*14+x*16+1],FIFO_1[256*14+x*16+1],FIFO_16[256*15+x*16+1],FIFO_15[256*15+x*16+1],FIFO_14[256*15+x*16+1],FIFO_13[256*15+x*16+1],FIFO_12[256*15+x*16+1],FIFO_11[256*15+x*16+1],FIFO_10[256*15+x*16+1],FIFO_9[256*15+x*16+1],FIFO_8[256*15+x*16+1],FIFO_7[256*15+x*16+1],FIFO_6[256*15+x*16+1],FIFO_5[256*15+x*16+1],FIFO_4[256*15+x*16+1],FIFO_3[256*15+x*16+1],FIFO_2[256*15+x*16+1],FIFO_1[256*15+x*16+1]}; 
                error_vector3 <= dec3 ^ {FIFO_16[256*0+x*16+2],FIFO_15[256*0+x*16+2],FIFO_14[256*0+x*16+2],FIFO_13[256*0+x*16+2],FIFO_12[256*0+x*16+2],FIFO_11[256*0+x*16+2],FIFO_10[256*0+x*16+2],FIFO_9[256*0+x*16+2],FIFO_8[256*0+x*16+2],FIFO_7[256*0+x*16+2],FIFO_6[256*0+x*16+2],FIFO_5[256*0+x*16+2],FIFO_4[256*0+x*16+2],FIFO_3[256*0+x*16+2],FIFO_2[256*0+x*16+2],FIFO_1[256*0+x*16+2],FIFO_16[256*1+x*16+2],FIFO_15[256*1+x*16+2],FIFO_14[256*1+x*16+2],FIFO_13[256*1+x*16+2],FIFO_12[256*1+x*16+2],FIFO_11[256*1+x*16+2],FIFO_10[256*1+x*16+2],FIFO_9[256*1+x*16+2],FIFO_8[256*1+x*16+2],FIFO_7[256*1+x*16+2],FIFO_6[256*1+x*16+2],FIFO_5[256*1+x*16+2],FIFO_4[256*1+x*16+2],FIFO_3[256*1+x*16+2],FIFO_2[256*1+x*16+2],FIFO_1[256*1+x*16+2],FIFO_16[256*2+x*16+2],FIFO_15[256*2+x*16+2],FIFO_14[256*2+x*16+2],FIFO_13[256*2+x*16+2],FIFO_12[256*2+x*16+2],FIFO_11[256*2+x*16+2],FIFO_10[256*2+x*16+2],FIFO_9[256*2+x*16+2],FIFO_8[256*2+x*16+2],FIFO_7[256*2+x*16+2],FIFO_6[256*2+x*16+2],FIFO_5[256*2+x*16+2],FIFO_4[256*2+x*16+2],FIFO_3[256*2+x*16+2],FIFO_2[256*2+x*16+2],FIFO_1[256*2+x*16+2],FIFO_16[256*3+x*16+2],FIFO_15[256*3+x*16+2],FIFO_14[256*3+x*16+2],FIFO_13[256*3+x*16+2],FIFO_12[256*3+x*16+2],FIFO_11[256*3+x*16+2],FIFO_10[256*3+x*16+2],FIFO_9[256*3+x*16+2],FIFO_8[256*3+x*16+2],FIFO_7[256*3+x*16+2],FIFO_6[256*3+x*16+2],FIFO_5[256*3+x*16+2],FIFO_4[256*3+x*16+2],FIFO_3[256*3+x*16+2],FIFO_2[256*3+x*16+2],FIFO_1[256*3+x*16+2],FIFO_16[256*4+x*16+2],FIFO_15[256*4+x*16+2],FIFO_14[256*4+x*16+2],FIFO_13[256*4+x*16+2],FIFO_12[256*4+x*16+2],FIFO_11[256*4+x*16+2],FIFO_10[256*4+x*16+2],FIFO_9[256*4+x*16+2],FIFO_8[256*4+x*16+2],FIFO_7[256*4+x*16+2],FIFO_6[256*4+x*16+2],FIFO_5[256*4+x*16+2],FIFO_4[256*4+x*16+2],FIFO_3[256*4+x*16+2],FIFO_2[256*4+x*16+2],FIFO_1[256*4+x*16+2],FIFO_16[256*5+x*16+2],FIFO_15[256*5+x*16+2],FIFO_14[256*5+x*16+2],FIFO_13[256*5+x*16+2],FIFO_12[256*5+x*16+2],FIFO_11[256*5+x*16+2],FIFO_10[256*5+x*16+2],FIFO_9[256*5+x*16+2],FIFO_8[256*5+x*16+2],FIFO_7[256*5+x*16+2],FIFO_6[256*5+x*16+2],FIFO_5[256*5+x*16+2],FIFO_4[256*5+x*16+2],FIFO_3[256*5+x*16+2],FIFO_2[256*5+x*16+2],FIFO_1[256*5+x*16+2],FIFO_16[256*6+x*16+2],FIFO_15[256*6+x*16+2],FIFO_14[256*6+x*16+2],FIFO_13[256*6+x*16+2],FIFO_12[256*6+x*16+2],FIFO_11[256*6+x*16+2],FIFO_10[256*6+x*16+2],FIFO_9[256*6+x*16+2],FIFO_8[256*6+x*16+2],FIFO_7[256*6+x*16+2],FIFO_6[256*6+x*16+2],FIFO_5[256*6+x*16+2],FIFO_4[256*6+x*16+2],FIFO_3[256*6+x*16+2],FIFO_2[256*6+x*16+2],FIFO_1[256*6+x*16+2],FIFO_16[256*7+x*16+2],FIFO_15[256*7+x*16+2],FIFO_14[256*7+x*16+2],FIFO_13[256*7+x*16+2],FIFO_12[256*7+x*16+2],FIFO_11[256*7+x*16+2],FIFO_10[256*7+x*16+2],FIFO_9[256*7+x*16+2],FIFO_8[256*7+x*16+2],FIFO_7[256*7+x*16+2],FIFO_6[256*7+x*16+2],FIFO_5[256*7+x*16+2],FIFO_4[256*7+x*16+2],FIFO_3[256*7+x*16+2],FIFO_2[256*7+x*16+2],FIFO_1[256*7+x*16+2],FIFO_16[256*8+x*16+2],FIFO_15[256*8+x*16+2],FIFO_14[256*8+x*16+2],FIFO_13[256*8+x*16+2],FIFO_12[256*8+x*16+2],FIFO_11[256*8+x*16+2],FIFO_10[256*8+x*16+2],FIFO_9[256*8+x*16+2],FIFO_8[256*8+x*16+2],FIFO_7[256*8+x*16+2],FIFO_6[256*8+x*16+2],FIFO_5[256*8+x*16+2],FIFO_4[256*8+x*16+2],FIFO_3[256*8+x*16+2],FIFO_2[256*8+x*16+2],FIFO_1[256*8+x*16+2],FIFO_16[256*9+x*16+2],FIFO_15[256*9+x*16+2],FIFO_14[256*9+x*16+2],FIFO_13[256*9+x*16+2],FIFO_12[256*9+x*16+2],FIFO_11[256*9+x*16+2],FIFO_10[256*9+x*16+2],FIFO_9[256*9+x*16+2],FIFO_8[256*9+x*16+2],FIFO_7[256*9+x*16+2],FIFO_6[256*9+x*16+2],FIFO_5[256*9+x*16+2],FIFO_4[256*9+x*16+2],FIFO_3[256*9+x*16+2],FIFO_2[256*9+x*16+2],FIFO_1[256*9+x*16+2],FIFO_16[256*10+x*16+2],FIFO_15[256*10+x*16+2],FIFO_14[256*10+x*16+2],FIFO_13[256*10+x*16+2],FIFO_12[256*10+x*16+2],FIFO_11[256*10+x*16+2],FIFO_10[256*10+x*16+2],FIFO_9[256*10+x*16+2],FIFO_8[256*10+x*16+2],FIFO_7[256*10+x*16+2],FIFO_6[256*10+x*16+2],FIFO_5[256*10+x*16+2],FIFO_4[256*10+x*16+2],FIFO_3[256*10+x*16+2],FIFO_2[256*10+x*16+2],FIFO_1[256*10+x*16+2],FIFO_16[256*11+x*16+2],FIFO_15[256*11+x*16+2],FIFO_14[256*11+x*16+2],FIFO_13[256*11+x*16+2],FIFO_12[256*11+x*16+2],FIFO_11[256*11+x*16+2],FIFO_10[256*11+x*16+2],FIFO_9[256*11+x*16+2],FIFO_8[256*11+x*16+2],FIFO_7[256*11+x*16+2],FIFO_6[256*11+x*16+2],FIFO_5[256*11+x*16+2],FIFO_4[256*11+x*16+2],FIFO_3[256*11+x*16+2],FIFO_2[256*11+x*16+2],FIFO_1[256*11+x*16+2],FIFO_16[256*12+x*16+2],FIFO_15[256*12+x*16+2],FIFO_14[256*12+x*16+2],FIFO_13[256*12+x*16+2],FIFO_12[256*12+x*16+2],FIFO_11[256*12+x*16+2],FIFO_10[256*12+x*16+2],FIFO_9[256*12+x*16+2],FIFO_8[256*12+x*16+2],FIFO_7[256*12+x*16+2],FIFO_6[256*12+x*16+2],FIFO_5[256*12+x*16+2],FIFO_4[256*12+x*16+2],FIFO_3[256*12+x*16+2],FIFO_2[256*12+x*16+2],FIFO_1[256*12+x*16+2],FIFO_16[256*13+x*16+2],FIFO_15[256*13+x*16+2],FIFO_14[256*13+x*16+2],FIFO_13[256*13+x*16+2],FIFO_12[256*13+x*16+2],FIFO_11[256*13+x*16+2],FIFO_10[256*13+x*16+2],FIFO_9[256*13+x*16+2],FIFO_8[256*13+x*16+2],FIFO_7[256*13+x*16+2],FIFO_6[256*13+x*16+2],FIFO_5[256*13+x*16+2],FIFO_4[256*13+x*16+2],FIFO_3[256*13+x*16+2],FIFO_2[256*13+x*16+2],FIFO_1[256*13+x*16+2],FIFO_16[256*14+x*16+2],FIFO_15[256*14+x*16+2],FIFO_14[256*14+x*16+2],FIFO_13[256*14+x*16+2],FIFO_12[256*14+x*16+2],FIFO_11[256*14+x*16+2],FIFO_10[256*14+x*16+2],FIFO_9[256*14+x*16+2],FIFO_8[256*14+x*16+2],FIFO_7[256*14+x*16+2],FIFO_6[256*14+x*16+2],FIFO_5[256*14+x*16+2],FIFO_4[256*14+x*16+2],FIFO_3[256*14+x*16+2],FIFO_2[256*14+x*16+2],FIFO_1[256*14+x*16+2],FIFO_16[256*15+x*16+2],FIFO_15[256*15+x*16+2],FIFO_14[256*15+x*16+2],FIFO_13[256*15+x*16+2],FIFO_12[256*15+x*16+2],FIFO_11[256*15+x*16+2],FIFO_10[256*15+x*16+2],FIFO_9[256*15+x*16+2],FIFO_8[256*15+x*16+2],FIFO_7[256*15+x*16+2],FIFO_6[256*15+x*16+2],FIFO_5[256*15+x*16+2],FIFO_4[256*15+x*16+2],FIFO_3[256*15+x*16+2],FIFO_2[256*15+x*16+2],FIFO_1[256*15+x*16+2]}; 
                error_vector4 <= dec4 ^ {FIFO_16[256*0+x*16+3],FIFO_15[256*0+x*16+3],FIFO_14[256*0+x*16+3],FIFO_13[256*0+x*16+3],FIFO_12[256*0+x*16+3],FIFO_11[256*0+x*16+3],FIFO_10[256*0+x*16+3],FIFO_9[256*0+x*16+3],FIFO_8[256*0+x*16+3],FIFO_7[256*0+x*16+3],FIFO_6[256*0+x*16+3],FIFO_5[256*0+x*16+3],FIFO_4[256*0+x*16+3],FIFO_3[256*0+x*16+3],FIFO_2[256*0+x*16+3],FIFO_1[256*0+x*16+3],FIFO_16[256*1+x*16+3],FIFO_15[256*1+x*16+3],FIFO_14[256*1+x*16+3],FIFO_13[256*1+x*16+3],FIFO_12[256*1+x*16+3],FIFO_11[256*1+x*16+3],FIFO_10[256*1+x*16+3],FIFO_9[256*1+x*16+3],FIFO_8[256*1+x*16+3],FIFO_7[256*1+x*16+3],FIFO_6[256*1+x*16+3],FIFO_5[256*1+x*16+3],FIFO_4[256*1+x*16+3],FIFO_3[256*1+x*16+3],FIFO_2[256*1+x*16+3],FIFO_1[256*1+x*16+3],FIFO_16[256*2+x*16+3],FIFO_15[256*2+x*16+3],FIFO_14[256*2+x*16+3],FIFO_13[256*2+x*16+3],FIFO_12[256*2+x*16+3],FIFO_11[256*2+x*16+3],FIFO_10[256*2+x*16+3],FIFO_9[256*2+x*16+3],FIFO_8[256*2+x*16+3],FIFO_7[256*2+x*16+3],FIFO_6[256*2+x*16+3],FIFO_5[256*2+x*16+3],FIFO_4[256*2+x*16+3],FIFO_3[256*2+x*16+3],FIFO_2[256*2+x*16+3],FIFO_1[256*2+x*16+3],FIFO_16[256*3+x*16+3],FIFO_15[256*3+x*16+3],FIFO_14[256*3+x*16+3],FIFO_13[256*3+x*16+3],FIFO_12[256*3+x*16+3],FIFO_11[256*3+x*16+3],FIFO_10[256*3+x*16+3],FIFO_9[256*3+x*16+3],FIFO_8[256*3+x*16+3],FIFO_7[256*3+x*16+3],FIFO_6[256*3+x*16+3],FIFO_5[256*3+x*16+3],FIFO_4[256*3+x*16+3],FIFO_3[256*3+x*16+3],FIFO_2[256*3+x*16+3],FIFO_1[256*3+x*16+3],FIFO_16[256*4+x*16+3],FIFO_15[256*4+x*16+3],FIFO_14[256*4+x*16+3],FIFO_13[256*4+x*16+3],FIFO_12[256*4+x*16+3],FIFO_11[256*4+x*16+3],FIFO_10[256*4+x*16+3],FIFO_9[256*4+x*16+3],FIFO_8[256*4+x*16+3],FIFO_7[256*4+x*16+3],FIFO_6[256*4+x*16+3],FIFO_5[256*4+x*16+3],FIFO_4[256*4+x*16+3],FIFO_3[256*4+x*16+3],FIFO_2[256*4+x*16+3],FIFO_1[256*4+x*16+3],FIFO_16[256*5+x*16+3],FIFO_15[256*5+x*16+3],FIFO_14[256*5+x*16+3],FIFO_13[256*5+x*16+3],FIFO_12[256*5+x*16+3],FIFO_11[256*5+x*16+3],FIFO_10[256*5+x*16+3],FIFO_9[256*5+x*16+3],FIFO_8[256*5+x*16+3],FIFO_7[256*5+x*16+3],FIFO_6[256*5+x*16+3],FIFO_5[256*5+x*16+3],FIFO_4[256*5+x*16+3],FIFO_3[256*5+x*16+3],FIFO_2[256*5+x*16+3],FIFO_1[256*5+x*16+3],FIFO_16[256*6+x*16+3],FIFO_15[256*6+x*16+3],FIFO_14[256*6+x*16+3],FIFO_13[256*6+x*16+3],FIFO_12[256*6+x*16+3],FIFO_11[256*6+x*16+3],FIFO_10[256*6+x*16+3],FIFO_9[256*6+x*16+3],FIFO_8[256*6+x*16+3],FIFO_7[256*6+x*16+3],FIFO_6[256*6+x*16+3],FIFO_5[256*6+x*16+3],FIFO_4[256*6+x*16+3],FIFO_3[256*6+x*16+3],FIFO_2[256*6+x*16+3],FIFO_1[256*6+x*16+3],FIFO_16[256*7+x*16+3],FIFO_15[256*7+x*16+3],FIFO_14[256*7+x*16+3],FIFO_13[256*7+x*16+3],FIFO_12[256*7+x*16+3],FIFO_11[256*7+x*16+3],FIFO_10[256*7+x*16+3],FIFO_9[256*7+x*16+3],FIFO_8[256*7+x*16+3],FIFO_7[256*7+x*16+3],FIFO_6[256*7+x*16+3],FIFO_5[256*7+x*16+3],FIFO_4[256*7+x*16+3],FIFO_3[256*7+x*16+3],FIFO_2[256*7+x*16+3],FIFO_1[256*7+x*16+3],FIFO_16[256*8+x*16+3],FIFO_15[256*8+x*16+3],FIFO_14[256*8+x*16+3],FIFO_13[256*8+x*16+3],FIFO_12[256*8+x*16+3],FIFO_11[256*8+x*16+3],FIFO_10[256*8+x*16+3],FIFO_9[256*8+x*16+3],FIFO_8[256*8+x*16+3],FIFO_7[256*8+x*16+3],FIFO_6[256*8+x*16+3],FIFO_5[256*8+x*16+3],FIFO_4[256*8+x*16+3],FIFO_3[256*8+x*16+3],FIFO_2[256*8+x*16+3],FIFO_1[256*8+x*16+3],FIFO_16[256*9+x*16+3],FIFO_15[256*9+x*16+3],FIFO_14[256*9+x*16+3],FIFO_13[256*9+x*16+3],FIFO_12[256*9+x*16+3],FIFO_11[256*9+x*16+3],FIFO_10[256*9+x*16+3],FIFO_9[256*9+x*16+3],FIFO_8[256*9+x*16+3],FIFO_7[256*9+x*16+3],FIFO_6[256*9+x*16+3],FIFO_5[256*9+x*16+3],FIFO_4[256*9+x*16+3],FIFO_3[256*9+x*16+3],FIFO_2[256*9+x*16+3],FIFO_1[256*9+x*16+3],FIFO_16[256*10+x*16+3],FIFO_15[256*10+x*16+3],FIFO_14[256*10+x*16+3],FIFO_13[256*10+x*16+3],FIFO_12[256*10+x*16+3],FIFO_11[256*10+x*16+3],FIFO_10[256*10+x*16+3],FIFO_9[256*10+x*16+3],FIFO_8[256*10+x*16+3],FIFO_7[256*10+x*16+3],FIFO_6[256*10+x*16+3],FIFO_5[256*10+x*16+3],FIFO_4[256*10+x*16+3],FIFO_3[256*10+x*16+3],FIFO_2[256*10+x*16+3],FIFO_1[256*10+x*16+3],FIFO_16[256*11+x*16+3],FIFO_15[256*11+x*16+3],FIFO_14[256*11+x*16+3],FIFO_13[256*11+x*16+3],FIFO_12[256*11+x*16+3],FIFO_11[256*11+x*16+3],FIFO_10[256*11+x*16+3],FIFO_9[256*11+x*16+3],FIFO_8[256*11+x*16+3],FIFO_7[256*11+x*16+3],FIFO_6[256*11+x*16+3],FIFO_5[256*11+x*16+3],FIFO_4[256*11+x*16+3],FIFO_3[256*11+x*16+3],FIFO_2[256*11+x*16+3],FIFO_1[256*11+x*16+3],FIFO_16[256*12+x*16+3],FIFO_15[256*12+x*16+3],FIFO_14[256*12+x*16+3],FIFO_13[256*12+x*16+3],FIFO_12[256*12+x*16+3],FIFO_11[256*12+x*16+3],FIFO_10[256*12+x*16+3],FIFO_9[256*12+x*16+3],FIFO_8[256*12+x*16+3],FIFO_7[256*12+x*16+3],FIFO_6[256*12+x*16+3],FIFO_5[256*12+x*16+3],FIFO_4[256*12+x*16+3],FIFO_3[256*12+x*16+3],FIFO_2[256*12+x*16+3],FIFO_1[256*12+x*16+3],FIFO_16[256*13+x*16+3],FIFO_15[256*13+x*16+3],FIFO_14[256*13+x*16+3],FIFO_13[256*13+x*16+3],FIFO_12[256*13+x*16+3],FIFO_11[256*13+x*16+3],FIFO_10[256*13+x*16+3],FIFO_9[256*13+x*16+3],FIFO_8[256*13+x*16+3],FIFO_7[256*13+x*16+3],FIFO_6[256*13+x*16+3],FIFO_5[256*13+x*16+3],FIFO_4[256*13+x*16+3],FIFO_3[256*13+x*16+3],FIFO_2[256*13+x*16+3],FIFO_1[256*13+x*16+3],FIFO_16[256*14+x*16+3],FIFO_15[256*14+x*16+3],FIFO_14[256*14+x*16+3],FIFO_13[256*14+x*16+3],FIFO_12[256*14+x*16+3],FIFO_11[256*14+x*16+3],FIFO_10[256*14+x*16+3],FIFO_9[256*14+x*16+3],FIFO_8[256*14+x*16+3],FIFO_7[256*14+x*16+3],FIFO_6[256*14+x*16+3],FIFO_5[256*14+x*16+3],FIFO_4[256*14+x*16+3],FIFO_3[256*14+x*16+3],FIFO_2[256*14+x*16+3],FIFO_1[256*14+x*16+3],FIFO_16[256*15+x*16+3],FIFO_15[256*15+x*16+3],FIFO_14[256*15+x*16+3],FIFO_13[256*15+x*16+3],FIFO_12[256*15+x*16+3],FIFO_11[256*15+x*16+3],FIFO_10[256*15+x*16+3],FIFO_9[256*15+x*16+3],FIFO_8[256*15+x*16+3],FIFO_7[256*15+x*16+3],FIFO_6[256*15+x*16+3],FIFO_5[256*15+x*16+3],FIFO_4[256*15+x*16+3],FIFO_3[256*15+x*16+3],FIFO_2[256*15+x*16+3],FIFO_1[256*15+x*16+3]}; 
                error_vector5 <= dec5 ^ {FIFO_16[256*0+x*16+4],FIFO_15[256*0+x*16+4],FIFO_14[256*0+x*16+4],FIFO_13[256*0+x*16+4],FIFO_12[256*0+x*16+4],FIFO_11[256*0+x*16+4],FIFO_10[256*0+x*16+4],FIFO_9[256*0+x*16+4],FIFO_8[256*0+x*16+4],FIFO_7[256*0+x*16+4],FIFO_6[256*0+x*16+4],FIFO_5[256*0+x*16+4],FIFO_4[256*0+x*16+4],FIFO_3[256*0+x*16+4],FIFO_2[256*0+x*16+4],FIFO_1[256*0+x*16+4],FIFO_16[256*1+x*16+4],FIFO_15[256*1+x*16+4],FIFO_14[256*1+x*16+4],FIFO_13[256*1+x*16+4],FIFO_12[256*1+x*16+4],FIFO_11[256*1+x*16+4],FIFO_10[256*1+x*16+4],FIFO_9[256*1+x*16+4],FIFO_8[256*1+x*16+4],FIFO_7[256*1+x*16+4],FIFO_6[256*1+x*16+4],FIFO_5[256*1+x*16+4],FIFO_4[256*1+x*16+4],FIFO_3[256*1+x*16+4],FIFO_2[256*1+x*16+4],FIFO_1[256*1+x*16+4],FIFO_16[256*2+x*16+4],FIFO_15[256*2+x*16+4],FIFO_14[256*2+x*16+4],FIFO_13[256*2+x*16+4],FIFO_12[256*2+x*16+4],FIFO_11[256*2+x*16+4],FIFO_10[256*2+x*16+4],FIFO_9[256*2+x*16+4],FIFO_8[256*2+x*16+4],FIFO_7[256*2+x*16+4],FIFO_6[256*2+x*16+4],FIFO_5[256*2+x*16+4],FIFO_4[256*2+x*16+4],FIFO_3[256*2+x*16+4],FIFO_2[256*2+x*16+4],FIFO_1[256*2+x*16+4],FIFO_16[256*3+x*16+4],FIFO_15[256*3+x*16+4],FIFO_14[256*3+x*16+4],FIFO_13[256*3+x*16+4],FIFO_12[256*3+x*16+4],FIFO_11[256*3+x*16+4],FIFO_10[256*3+x*16+4],FIFO_9[256*3+x*16+4],FIFO_8[256*3+x*16+4],FIFO_7[256*3+x*16+4],FIFO_6[256*3+x*16+4],FIFO_5[256*3+x*16+4],FIFO_4[256*3+x*16+4],FIFO_3[256*3+x*16+4],FIFO_2[256*3+x*16+4],FIFO_1[256*3+x*16+4],FIFO_16[256*4+x*16+4],FIFO_15[256*4+x*16+4],FIFO_14[256*4+x*16+4],FIFO_13[256*4+x*16+4],FIFO_12[256*4+x*16+4],FIFO_11[256*4+x*16+4],FIFO_10[256*4+x*16+4],FIFO_9[256*4+x*16+4],FIFO_8[256*4+x*16+4],FIFO_7[256*4+x*16+4],FIFO_6[256*4+x*16+4],FIFO_5[256*4+x*16+4],FIFO_4[256*4+x*16+4],FIFO_3[256*4+x*16+4],FIFO_2[256*4+x*16+4],FIFO_1[256*4+x*16+4],FIFO_16[256*5+x*16+4],FIFO_15[256*5+x*16+4],FIFO_14[256*5+x*16+4],FIFO_13[256*5+x*16+4],FIFO_12[256*5+x*16+4],FIFO_11[256*5+x*16+4],FIFO_10[256*5+x*16+4],FIFO_9[256*5+x*16+4],FIFO_8[256*5+x*16+4],FIFO_7[256*5+x*16+4],FIFO_6[256*5+x*16+4],FIFO_5[256*5+x*16+4],FIFO_4[256*5+x*16+4],FIFO_3[256*5+x*16+4],FIFO_2[256*5+x*16+4],FIFO_1[256*5+x*16+4],FIFO_16[256*6+x*16+4],FIFO_15[256*6+x*16+4],FIFO_14[256*6+x*16+4],FIFO_13[256*6+x*16+4],FIFO_12[256*6+x*16+4],FIFO_11[256*6+x*16+4],FIFO_10[256*6+x*16+4],FIFO_9[256*6+x*16+4],FIFO_8[256*6+x*16+4],FIFO_7[256*6+x*16+4],FIFO_6[256*6+x*16+4],FIFO_5[256*6+x*16+4],FIFO_4[256*6+x*16+4],FIFO_3[256*6+x*16+4],FIFO_2[256*6+x*16+4],FIFO_1[256*6+x*16+4],FIFO_16[256*7+x*16+4],FIFO_15[256*7+x*16+4],FIFO_14[256*7+x*16+4],FIFO_13[256*7+x*16+4],FIFO_12[256*7+x*16+4],FIFO_11[256*7+x*16+4],FIFO_10[256*7+x*16+4],FIFO_9[256*7+x*16+4],FIFO_8[256*7+x*16+4],FIFO_7[256*7+x*16+4],FIFO_6[256*7+x*16+4],FIFO_5[256*7+x*16+4],FIFO_4[256*7+x*16+4],FIFO_3[256*7+x*16+4],FIFO_2[256*7+x*16+4],FIFO_1[256*7+x*16+4],FIFO_16[256*8+x*16+4],FIFO_15[256*8+x*16+4],FIFO_14[256*8+x*16+4],FIFO_13[256*8+x*16+4],FIFO_12[256*8+x*16+4],FIFO_11[256*8+x*16+4],FIFO_10[256*8+x*16+4],FIFO_9[256*8+x*16+4],FIFO_8[256*8+x*16+4],FIFO_7[256*8+x*16+4],FIFO_6[256*8+x*16+4],FIFO_5[256*8+x*16+4],FIFO_4[256*8+x*16+4],FIFO_3[256*8+x*16+4],FIFO_2[256*8+x*16+4],FIFO_1[256*8+x*16+4],FIFO_16[256*9+x*16+4],FIFO_15[256*9+x*16+4],FIFO_14[256*9+x*16+4],FIFO_13[256*9+x*16+4],FIFO_12[256*9+x*16+4],FIFO_11[256*9+x*16+4],FIFO_10[256*9+x*16+4],FIFO_9[256*9+x*16+4],FIFO_8[256*9+x*16+4],FIFO_7[256*9+x*16+4],FIFO_6[256*9+x*16+4],FIFO_5[256*9+x*16+4],FIFO_4[256*9+x*16+4],FIFO_3[256*9+x*16+4],FIFO_2[256*9+x*16+4],FIFO_1[256*9+x*16+4],FIFO_16[256*10+x*16+4],FIFO_15[256*10+x*16+4],FIFO_14[256*10+x*16+4],FIFO_13[256*10+x*16+4],FIFO_12[256*10+x*16+4],FIFO_11[256*10+x*16+4],FIFO_10[256*10+x*16+4],FIFO_9[256*10+x*16+4],FIFO_8[256*10+x*16+4],FIFO_7[256*10+x*16+4],FIFO_6[256*10+x*16+4],FIFO_5[256*10+x*16+4],FIFO_4[256*10+x*16+4],FIFO_3[256*10+x*16+4],FIFO_2[256*10+x*16+4],FIFO_1[256*10+x*16+4],FIFO_16[256*11+x*16+4],FIFO_15[256*11+x*16+4],FIFO_14[256*11+x*16+4],FIFO_13[256*11+x*16+4],FIFO_12[256*11+x*16+4],FIFO_11[256*11+x*16+4],FIFO_10[256*11+x*16+4],FIFO_9[256*11+x*16+4],FIFO_8[256*11+x*16+4],FIFO_7[256*11+x*16+4],FIFO_6[256*11+x*16+4],FIFO_5[256*11+x*16+4],FIFO_4[256*11+x*16+4],FIFO_3[256*11+x*16+4],FIFO_2[256*11+x*16+4],FIFO_1[256*11+x*16+4],FIFO_16[256*12+x*16+4],FIFO_15[256*12+x*16+4],FIFO_14[256*12+x*16+4],FIFO_13[256*12+x*16+4],FIFO_12[256*12+x*16+4],FIFO_11[256*12+x*16+4],FIFO_10[256*12+x*16+4],FIFO_9[256*12+x*16+4],FIFO_8[256*12+x*16+4],FIFO_7[256*12+x*16+4],FIFO_6[256*12+x*16+4],FIFO_5[256*12+x*16+4],FIFO_4[256*12+x*16+4],FIFO_3[256*12+x*16+4],FIFO_2[256*12+x*16+4],FIFO_1[256*12+x*16+4],FIFO_16[256*13+x*16+4],FIFO_15[256*13+x*16+4],FIFO_14[256*13+x*16+4],FIFO_13[256*13+x*16+4],FIFO_12[256*13+x*16+4],FIFO_11[256*13+x*16+4],FIFO_10[256*13+x*16+4],FIFO_9[256*13+x*16+4],FIFO_8[256*13+x*16+4],FIFO_7[256*13+x*16+4],FIFO_6[256*13+x*16+4],FIFO_5[256*13+x*16+4],FIFO_4[256*13+x*16+4],FIFO_3[256*13+x*16+4],FIFO_2[256*13+x*16+4],FIFO_1[256*13+x*16+4],FIFO_16[256*14+x*16+4],FIFO_15[256*14+x*16+4],FIFO_14[256*14+x*16+4],FIFO_13[256*14+x*16+4],FIFO_12[256*14+x*16+4],FIFO_11[256*14+x*16+4],FIFO_10[256*14+x*16+4],FIFO_9[256*14+x*16+4],FIFO_8[256*14+x*16+4],FIFO_7[256*14+x*16+4],FIFO_6[256*14+x*16+4],FIFO_5[256*14+x*16+4],FIFO_4[256*14+x*16+4],FIFO_3[256*14+x*16+4],FIFO_2[256*14+x*16+4],FIFO_1[256*14+x*16+4],FIFO_16[256*15+x*16+4],FIFO_15[256*15+x*16+4],FIFO_14[256*15+x*16+4],FIFO_13[256*15+x*16+4],FIFO_12[256*15+x*16+4],FIFO_11[256*15+x*16+4],FIFO_10[256*15+x*16+4],FIFO_9[256*15+x*16+4],FIFO_8[256*15+x*16+4],FIFO_7[256*15+x*16+4],FIFO_6[256*15+x*16+4],FIFO_5[256*15+x*16+4],FIFO_4[256*15+x*16+4],FIFO_3[256*15+x*16+4],FIFO_2[256*15+x*16+4],FIFO_1[256*15+x*16+4]}; 
                error_vector6 <= dec6 ^ {FIFO_16[256*0+x*16+5],FIFO_15[256*0+x*16+5],FIFO_14[256*0+x*16+5],FIFO_13[256*0+x*16+5],FIFO_12[256*0+x*16+5],FIFO_11[256*0+x*16+5],FIFO_10[256*0+x*16+5],FIFO_9[256*0+x*16+5],FIFO_8[256*0+x*16+5],FIFO_7[256*0+x*16+5],FIFO_6[256*0+x*16+5],FIFO_5[256*0+x*16+5],FIFO_4[256*0+x*16+5],FIFO_3[256*0+x*16+5],FIFO_2[256*0+x*16+5],FIFO_1[256*0+x*16+5],FIFO_16[256*1+x*16+5],FIFO_15[256*1+x*16+5],FIFO_14[256*1+x*16+5],FIFO_13[256*1+x*16+5],FIFO_12[256*1+x*16+5],FIFO_11[256*1+x*16+5],FIFO_10[256*1+x*16+5],FIFO_9[256*1+x*16+5],FIFO_8[256*1+x*16+5],FIFO_7[256*1+x*16+5],FIFO_6[256*1+x*16+5],FIFO_5[256*1+x*16+5],FIFO_4[256*1+x*16+5],FIFO_3[256*1+x*16+5],FIFO_2[256*1+x*16+5],FIFO_1[256*1+x*16+5],FIFO_16[256*2+x*16+5],FIFO_15[256*2+x*16+5],FIFO_14[256*2+x*16+5],FIFO_13[256*2+x*16+5],FIFO_12[256*2+x*16+5],FIFO_11[256*2+x*16+5],FIFO_10[256*2+x*16+5],FIFO_9[256*2+x*16+5],FIFO_8[256*2+x*16+5],FIFO_7[256*2+x*16+5],FIFO_6[256*2+x*16+5],FIFO_5[256*2+x*16+5],FIFO_4[256*2+x*16+5],FIFO_3[256*2+x*16+5],FIFO_2[256*2+x*16+5],FIFO_1[256*2+x*16+5],FIFO_16[256*3+x*16+5],FIFO_15[256*3+x*16+5],FIFO_14[256*3+x*16+5],FIFO_13[256*3+x*16+5],FIFO_12[256*3+x*16+5],FIFO_11[256*3+x*16+5],FIFO_10[256*3+x*16+5],FIFO_9[256*3+x*16+5],FIFO_8[256*3+x*16+5],FIFO_7[256*3+x*16+5],FIFO_6[256*3+x*16+5],FIFO_5[256*3+x*16+5],FIFO_4[256*3+x*16+5],FIFO_3[256*3+x*16+5],FIFO_2[256*3+x*16+5],FIFO_1[256*3+x*16+5],FIFO_16[256*4+x*16+5],FIFO_15[256*4+x*16+5],FIFO_14[256*4+x*16+5],FIFO_13[256*4+x*16+5],FIFO_12[256*4+x*16+5],FIFO_11[256*4+x*16+5],FIFO_10[256*4+x*16+5],FIFO_9[256*4+x*16+5],FIFO_8[256*4+x*16+5],FIFO_7[256*4+x*16+5],FIFO_6[256*4+x*16+5],FIFO_5[256*4+x*16+5],FIFO_4[256*4+x*16+5],FIFO_3[256*4+x*16+5],FIFO_2[256*4+x*16+5],FIFO_1[256*4+x*16+5],FIFO_16[256*5+x*16+5],FIFO_15[256*5+x*16+5],FIFO_14[256*5+x*16+5],FIFO_13[256*5+x*16+5],FIFO_12[256*5+x*16+5],FIFO_11[256*5+x*16+5],FIFO_10[256*5+x*16+5],FIFO_9[256*5+x*16+5],FIFO_8[256*5+x*16+5],FIFO_7[256*5+x*16+5],FIFO_6[256*5+x*16+5],FIFO_5[256*5+x*16+5],FIFO_4[256*5+x*16+5],FIFO_3[256*5+x*16+5],FIFO_2[256*5+x*16+5],FIFO_1[256*5+x*16+5],FIFO_16[256*6+x*16+5],FIFO_15[256*6+x*16+5],FIFO_14[256*6+x*16+5],FIFO_13[256*6+x*16+5],FIFO_12[256*6+x*16+5],FIFO_11[256*6+x*16+5],FIFO_10[256*6+x*16+5],FIFO_9[256*6+x*16+5],FIFO_8[256*6+x*16+5],FIFO_7[256*6+x*16+5],FIFO_6[256*6+x*16+5],FIFO_5[256*6+x*16+5],FIFO_4[256*6+x*16+5],FIFO_3[256*6+x*16+5],FIFO_2[256*6+x*16+5],FIFO_1[256*6+x*16+5],FIFO_16[256*7+x*16+5],FIFO_15[256*7+x*16+5],FIFO_14[256*7+x*16+5],FIFO_13[256*7+x*16+5],FIFO_12[256*7+x*16+5],FIFO_11[256*7+x*16+5],FIFO_10[256*7+x*16+5],FIFO_9[256*7+x*16+5],FIFO_8[256*7+x*16+5],FIFO_7[256*7+x*16+5],FIFO_6[256*7+x*16+5],FIFO_5[256*7+x*16+5],FIFO_4[256*7+x*16+5],FIFO_3[256*7+x*16+5],FIFO_2[256*7+x*16+5],FIFO_1[256*7+x*16+5],FIFO_16[256*8+x*16+5],FIFO_15[256*8+x*16+5],FIFO_14[256*8+x*16+5],FIFO_13[256*8+x*16+5],FIFO_12[256*8+x*16+5],FIFO_11[256*8+x*16+5],FIFO_10[256*8+x*16+5],FIFO_9[256*8+x*16+5],FIFO_8[256*8+x*16+5],FIFO_7[256*8+x*16+5],FIFO_6[256*8+x*16+5],FIFO_5[256*8+x*16+5],FIFO_4[256*8+x*16+5],FIFO_3[256*8+x*16+5],FIFO_2[256*8+x*16+5],FIFO_1[256*8+x*16+5],FIFO_16[256*9+x*16+5],FIFO_15[256*9+x*16+5],FIFO_14[256*9+x*16+5],FIFO_13[256*9+x*16+5],FIFO_12[256*9+x*16+5],FIFO_11[256*9+x*16+5],FIFO_10[256*9+x*16+5],FIFO_9[256*9+x*16+5],FIFO_8[256*9+x*16+5],FIFO_7[256*9+x*16+5],FIFO_6[256*9+x*16+5],FIFO_5[256*9+x*16+5],FIFO_4[256*9+x*16+5],FIFO_3[256*9+x*16+5],FIFO_2[256*9+x*16+5],FIFO_1[256*9+x*16+5],FIFO_16[256*10+x*16+5],FIFO_15[256*10+x*16+5],FIFO_14[256*10+x*16+5],FIFO_13[256*10+x*16+5],FIFO_12[256*10+x*16+5],FIFO_11[256*10+x*16+5],FIFO_10[256*10+x*16+5],FIFO_9[256*10+x*16+5],FIFO_8[256*10+x*16+5],FIFO_7[256*10+x*16+5],FIFO_6[256*10+x*16+5],FIFO_5[256*10+x*16+5],FIFO_4[256*10+x*16+5],FIFO_3[256*10+x*16+5],FIFO_2[256*10+x*16+5],FIFO_1[256*10+x*16+5],FIFO_16[256*11+x*16+5],FIFO_15[256*11+x*16+5],FIFO_14[256*11+x*16+5],FIFO_13[256*11+x*16+5],FIFO_12[256*11+x*16+5],FIFO_11[256*11+x*16+5],FIFO_10[256*11+x*16+5],FIFO_9[256*11+x*16+5],FIFO_8[256*11+x*16+5],FIFO_7[256*11+x*16+5],FIFO_6[256*11+x*16+5],FIFO_5[256*11+x*16+5],FIFO_4[256*11+x*16+5],FIFO_3[256*11+x*16+5],FIFO_2[256*11+x*16+5],FIFO_1[256*11+x*16+5],FIFO_16[256*12+x*16+5],FIFO_15[256*12+x*16+5],FIFO_14[256*12+x*16+5],FIFO_13[256*12+x*16+5],FIFO_12[256*12+x*16+5],FIFO_11[256*12+x*16+5],FIFO_10[256*12+x*16+5],FIFO_9[256*12+x*16+5],FIFO_8[256*12+x*16+5],FIFO_7[256*12+x*16+5],FIFO_6[256*12+x*16+5],FIFO_5[256*12+x*16+5],FIFO_4[256*12+x*16+5],FIFO_3[256*12+x*16+5],FIFO_2[256*12+x*16+5],FIFO_1[256*12+x*16+5],FIFO_16[256*13+x*16+5],FIFO_15[256*13+x*16+5],FIFO_14[256*13+x*16+5],FIFO_13[256*13+x*16+5],FIFO_12[256*13+x*16+5],FIFO_11[256*13+x*16+5],FIFO_10[256*13+x*16+5],FIFO_9[256*13+x*16+5],FIFO_8[256*13+x*16+5],FIFO_7[256*13+x*16+5],FIFO_6[256*13+x*16+5],FIFO_5[256*13+x*16+5],FIFO_4[256*13+x*16+5],FIFO_3[256*13+x*16+5],FIFO_2[256*13+x*16+5],FIFO_1[256*13+x*16+5],FIFO_16[256*14+x*16+5],FIFO_15[256*14+x*16+5],FIFO_14[256*14+x*16+5],FIFO_13[256*14+x*16+5],FIFO_12[256*14+x*16+5],FIFO_11[256*14+x*16+5],FIFO_10[256*14+x*16+5],FIFO_9[256*14+x*16+5],FIFO_8[256*14+x*16+5],FIFO_7[256*14+x*16+5],FIFO_6[256*14+x*16+5],FIFO_5[256*14+x*16+5],FIFO_4[256*14+x*16+5],FIFO_3[256*14+x*16+5],FIFO_2[256*14+x*16+5],FIFO_1[256*14+x*16+5],FIFO_16[256*15+x*16+5],FIFO_15[256*15+x*16+5],FIFO_14[256*15+x*16+5],FIFO_13[256*15+x*16+5],FIFO_12[256*15+x*16+5],FIFO_11[256*15+x*16+5],FIFO_10[256*15+x*16+5],FIFO_9[256*15+x*16+5],FIFO_8[256*15+x*16+5],FIFO_7[256*15+x*16+5],FIFO_6[256*15+x*16+5],FIFO_5[256*15+x*16+5],FIFO_4[256*15+x*16+5],FIFO_3[256*15+x*16+5],FIFO_2[256*15+x*16+5],FIFO_1[256*15+x*16+5]}; 
                error_vector7 <= dec7 ^ {FIFO_16[256*0+x*16+6],FIFO_15[256*0+x*16+6],FIFO_14[256*0+x*16+6],FIFO_13[256*0+x*16+6],FIFO_12[256*0+x*16+6],FIFO_11[256*0+x*16+6],FIFO_10[256*0+x*16+6],FIFO_9[256*0+x*16+6],FIFO_8[256*0+x*16+6],FIFO_7[256*0+x*16+6],FIFO_6[256*0+x*16+6],FIFO_5[256*0+x*16+6],FIFO_4[256*0+x*16+6],FIFO_3[256*0+x*16+6],FIFO_2[256*0+x*16+6],FIFO_1[256*0+x*16+6],FIFO_16[256*1+x*16+6],FIFO_15[256*1+x*16+6],FIFO_14[256*1+x*16+6],FIFO_13[256*1+x*16+6],FIFO_12[256*1+x*16+6],FIFO_11[256*1+x*16+6],FIFO_10[256*1+x*16+6],FIFO_9[256*1+x*16+6],FIFO_8[256*1+x*16+6],FIFO_7[256*1+x*16+6],FIFO_6[256*1+x*16+6],FIFO_5[256*1+x*16+6],FIFO_4[256*1+x*16+6],FIFO_3[256*1+x*16+6],FIFO_2[256*1+x*16+6],FIFO_1[256*1+x*16+6],FIFO_16[256*2+x*16+6],FIFO_15[256*2+x*16+6],FIFO_14[256*2+x*16+6],FIFO_13[256*2+x*16+6],FIFO_12[256*2+x*16+6],FIFO_11[256*2+x*16+6],FIFO_10[256*2+x*16+6],FIFO_9[256*2+x*16+6],FIFO_8[256*2+x*16+6],FIFO_7[256*2+x*16+6],FIFO_6[256*2+x*16+6],FIFO_5[256*2+x*16+6],FIFO_4[256*2+x*16+6],FIFO_3[256*2+x*16+6],FIFO_2[256*2+x*16+6],FIFO_1[256*2+x*16+6],FIFO_16[256*3+x*16+6],FIFO_15[256*3+x*16+6],FIFO_14[256*3+x*16+6],FIFO_13[256*3+x*16+6],FIFO_12[256*3+x*16+6],FIFO_11[256*3+x*16+6],FIFO_10[256*3+x*16+6],FIFO_9[256*3+x*16+6],FIFO_8[256*3+x*16+6],FIFO_7[256*3+x*16+6],FIFO_6[256*3+x*16+6],FIFO_5[256*3+x*16+6],FIFO_4[256*3+x*16+6],FIFO_3[256*3+x*16+6],FIFO_2[256*3+x*16+6],FIFO_1[256*3+x*16+6],FIFO_16[256*4+x*16+6],FIFO_15[256*4+x*16+6],FIFO_14[256*4+x*16+6],FIFO_13[256*4+x*16+6],FIFO_12[256*4+x*16+6],FIFO_11[256*4+x*16+6],FIFO_10[256*4+x*16+6],FIFO_9[256*4+x*16+6],FIFO_8[256*4+x*16+6],FIFO_7[256*4+x*16+6],FIFO_6[256*4+x*16+6],FIFO_5[256*4+x*16+6],FIFO_4[256*4+x*16+6],FIFO_3[256*4+x*16+6],FIFO_2[256*4+x*16+6],FIFO_1[256*4+x*16+6],FIFO_16[256*5+x*16+6],FIFO_15[256*5+x*16+6],FIFO_14[256*5+x*16+6],FIFO_13[256*5+x*16+6],FIFO_12[256*5+x*16+6],FIFO_11[256*5+x*16+6],FIFO_10[256*5+x*16+6],FIFO_9[256*5+x*16+6],FIFO_8[256*5+x*16+6],FIFO_7[256*5+x*16+6],FIFO_6[256*5+x*16+6],FIFO_5[256*5+x*16+6],FIFO_4[256*5+x*16+6],FIFO_3[256*5+x*16+6],FIFO_2[256*5+x*16+6],FIFO_1[256*5+x*16+6],FIFO_16[256*6+x*16+6],FIFO_15[256*6+x*16+6],FIFO_14[256*6+x*16+6],FIFO_13[256*6+x*16+6],FIFO_12[256*6+x*16+6],FIFO_11[256*6+x*16+6],FIFO_10[256*6+x*16+6],FIFO_9[256*6+x*16+6],FIFO_8[256*6+x*16+6],FIFO_7[256*6+x*16+6],FIFO_6[256*6+x*16+6],FIFO_5[256*6+x*16+6],FIFO_4[256*6+x*16+6],FIFO_3[256*6+x*16+6],FIFO_2[256*6+x*16+6],FIFO_1[256*6+x*16+6],FIFO_16[256*7+x*16+6],FIFO_15[256*7+x*16+6],FIFO_14[256*7+x*16+6],FIFO_13[256*7+x*16+6],FIFO_12[256*7+x*16+6],FIFO_11[256*7+x*16+6],FIFO_10[256*7+x*16+6],FIFO_9[256*7+x*16+6],FIFO_8[256*7+x*16+6],FIFO_7[256*7+x*16+6],FIFO_6[256*7+x*16+6],FIFO_5[256*7+x*16+6],FIFO_4[256*7+x*16+6],FIFO_3[256*7+x*16+6],FIFO_2[256*7+x*16+6],FIFO_1[256*7+x*16+6],FIFO_16[256*8+x*16+6],FIFO_15[256*8+x*16+6],FIFO_14[256*8+x*16+6],FIFO_13[256*8+x*16+6],FIFO_12[256*8+x*16+6],FIFO_11[256*8+x*16+6],FIFO_10[256*8+x*16+6],FIFO_9[256*8+x*16+6],FIFO_8[256*8+x*16+6],FIFO_7[256*8+x*16+6],FIFO_6[256*8+x*16+6],FIFO_5[256*8+x*16+6],FIFO_4[256*8+x*16+6],FIFO_3[256*8+x*16+6],FIFO_2[256*8+x*16+6],FIFO_1[256*8+x*16+6],FIFO_16[256*9+x*16+6],FIFO_15[256*9+x*16+6],FIFO_14[256*9+x*16+6],FIFO_13[256*9+x*16+6],FIFO_12[256*9+x*16+6],FIFO_11[256*9+x*16+6],FIFO_10[256*9+x*16+6],FIFO_9[256*9+x*16+6],FIFO_8[256*9+x*16+6],FIFO_7[256*9+x*16+6],FIFO_6[256*9+x*16+6],FIFO_5[256*9+x*16+6],FIFO_4[256*9+x*16+6],FIFO_3[256*9+x*16+6],FIFO_2[256*9+x*16+6],FIFO_1[256*9+x*16+6],FIFO_16[256*10+x*16+6],FIFO_15[256*10+x*16+6],FIFO_14[256*10+x*16+6],FIFO_13[256*10+x*16+6],FIFO_12[256*10+x*16+6],FIFO_11[256*10+x*16+6],FIFO_10[256*10+x*16+6],FIFO_9[256*10+x*16+6],FIFO_8[256*10+x*16+6],FIFO_7[256*10+x*16+6],FIFO_6[256*10+x*16+6],FIFO_5[256*10+x*16+6],FIFO_4[256*10+x*16+6],FIFO_3[256*10+x*16+6],FIFO_2[256*10+x*16+6],FIFO_1[256*10+x*16+6],FIFO_16[256*11+x*16+6],FIFO_15[256*11+x*16+6],FIFO_14[256*11+x*16+6],FIFO_13[256*11+x*16+6],FIFO_12[256*11+x*16+6],FIFO_11[256*11+x*16+6],FIFO_10[256*11+x*16+6],FIFO_9[256*11+x*16+6],FIFO_8[256*11+x*16+6],FIFO_7[256*11+x*16+6],FIFO_6[256*11+x*16+6],FIFO_5[256*11+x*16+6],FIFO_4[256*11+x*16+6],FIFO_3[256*11+x*16+6],FIFO_2[256*11+x*16+6],FIFO_1[256*11+x*16+6],FIFO_16[256*12+x*16+6],FIFO_15[256*12+x*16+6],FIFO_14[256*12+x*16+6],FIFO_13[256*12+x*16+6],FIFO_12[256*12+x*16+6],FIFO_11[256*12+x*16+6],FIFO_10[256*12+x*16+6],FIFO_9[256*12+x*16+6],FIFO_8[256*12+x*16+6],FIFO_7[256*12+x*16+6],FIFO_6[256*12+x*16+6],FIFO_5[256*12+x*16+6],FIFO_4[256*12+x*16+6],FIFO_3[256*12+x*16+6],FIFO_2[256*12+x*16+6],FIFO_1[256*12+x*16+6],FIFO_16[256*13+x*16+6],FIFO_15[256*13+x*16+6],FIFO_14[256*13+x*16+6],FIFO_13[256*13+x*16+6],FIFO_12[256*13+x*16+6],FIFO_11[256*13+x*16+6],FIFO_10[256*13+x*16+6],FIFO_9[256*13+x*16+6],FIFO_8[256*13+x*16+6],FIFO_7[256*13+x*16+6],FIFO_6[256*13+x*16+6],FIFO_5[256*13+x*16+6],FIFO_4[256*13+x*16+6],FIFO_3[256*13+x*16+6],FIFO_2[256*13+x*16+6],FIFO_1[256*13+x*16+6],FIFO_16[256*14+x*16+6],FIFO_15[256*14+x*16+6],FIFO_14[256*14+x*16+6],FIFO_13[256*14+x*16+6],FIFO_12[256*14+x*16+6],FIFO_11[256*14+x*16+6],FIFO_10[256*14+x*16+6],FIFO_9[256*14+x*16+6],FIFO_8[256*14+x*16+6],FIFO_7[256*14+x*16+6],FIFO_6[256*14+x*16+6],FIFO_5[256*14+x*16+6],FIFO_4[256*14+x*16+6],FIFO_3[256*14+x*16+6],FIFO_2[256*14+x*16+6],FIFO_1[256*14+x*16+6],FIFO_16[256*15+x*16+6],FIFO_15[256*15+x*16+6],FIFO_14[256*15+x*16+6],FIFO_13[256*15+x*16+6],FIFO_12[256*15+x*16+6],FIFO_11[256*15+x*16+6],FIFO_10[256*15+x*16+6],FIFO_9[256*15+x*16+6],FIFO_8[256*15+x*16+6],FIFO_7[256*15+x*16+6],FIFO_6[256*15+x*16+6],FIFO_5[256*15+x*16+6],FIFO_4[256*15+x*16+6],FIFO_3[256*15+x*16+6],FIFO_2[256*15+x*16+6],FIFO_1[256*15+x*16+6]}; 
                error_vector8 <= dec8 ^ {FIFO_16[256*0+x*16+7],FIFO_15[256*0+x*16+7],FIFO_14[256*0+x*16+7],FIFO_13[256*0+x*16+7],FIFO_12[256*0+x*16+7],FIFO_11[256*0+x*16+7],FIFO_10[256*0+x*16+7],FIFO_9[256*0+x*16+7],FIFO_8[256*0+x*16+7],FIFO_7[256*0+x*16+7],FIFO_6[256*0+x*16+7],FIFO_5[256*0+x*16+7],FIFO_4[256*0+x*16+7],FIFO_3[256*0+x*16+7],FIFO_2[256*0+x*16+7],FIFO_1[256*0+x*16+7],FIFO_16[256*1+x*16+7],FIFO_15[256*1+x*16+7],FIFO_14[256*1+x*16+7],FIFO_13[256*1+x*16+7],FIFO_12[256*1+x*16+7],FIFO_11[256*1+x*16+7],FIFO_10[256*1+x*16+7],FIFO_9[256*1+x*16+7],FIFO_8[256*1+x*16+7],FIFO_7[256*1+x*16+7],FIFO_6[256*1+x*16+7],FIFO_5[256*1+x*16+7],FIFO_4[256*1+x*16+7],FIFO_3[256*1+x*16+7],FIFO_2[256*1+x*16+7],FIFO_1[256*1+x*16+7],FIFO_16[256*2+x*16+7],FIFO_15[256*2+x*16+7],FIFO_14[256*2+x*16+7],FIFO_13[256*2+x*16+7],FIFO_12[256*2+x*16+7],FIFO_11[256*2+x*16+7],FIFO_10[256*2+x*16+7],FIFO_9[256*2+x*16+7],FIFO_8[256*2+x*16+7],FIFO_7[256*2+x*16+7],FIFO_6[256*2+x*16+7],FIFO_5[256*2+x*16+7],FIFO_4[256*2+x*16+7],FIFO_3[256*2+x*16+7],FIFO_2[256*2+x*16+7],FIFO_1[256*2+x*16+7],FIFO_16[256*3+x*16+7],FIFO_15[256*3+x*16+7],FIFO_14[256*3+x*16+7],FIFO_13[256*3+x*16+7],FIFO_12[256*3+x*16+7],FIFO_11[256*3+x*16+7],FIFO_10[256*3+x*16+7],FIFO_9[256*3+x*16+7],FIFO_8[256*3+x*16+7],FIFO_7[256*3+x*16+7],FIFO_6[256*3+x*16+7],FIFO_5[256*3+x*16+7],FIFO_4[256*3+x*16+7],FIFO_3[256*3+x*16+7],FIFO_2[256*3+x*16+7],FIFO_1[256*3+x*16+7],FIFO_16[256*4+x*16+7],FIFO_15[256*4+x*16+7],FIFO_14[256*4+x*16+7],FIFO_13[256*4+x*16+7],FIFO_12[256*4+x*16+7],FIFO_11[256*4+x*16+7],FIFO_10[256*4+x*16+7],FIFO_9[256*4+x*16+7],FIFO_8[256*4+x*16+7],FIFO_7[256*4+x*16+7],FIFO_6[256*4+x*16+7],FIFO_5[256*4+x*16+7],FIFO_4[256*4+x*16+7],FIFO_3[256*4+x*16+7],FIFO_2[256*4+x*16+7],FIFO_1[256*4+x*16+7],FIFO_16[256*5+x*16+7],FIFO_15[256*5+x*16+7],FIFO_14[256*5+x*16+7],FIFO_13[256*5+x*16+7],FIFO_12[256*5+x*16+7],FIFO_11[256*5+x*16+7],FIFO_10[256*5+x*16+7],FIFO_9[256*5+x*16+7],FIFO_8[256*5+x*16+7],FIFO_7[256*5+x*16+7],FIFO_6[256*5+x*16+7],FIFO_5[256*5+x*16+7],FIFO_4[256*5+x*16+7],FIFO_3[256*5+x*16+7],FIFO_2[256*5+x*16+7],FIFO_1[256*5+x*16+7],FIFO_16[256*6+x*16+7],FIFO_15[256*6+x*16+7],FIFO_14[256*6+x*16+7],FIFO_13[256*6+x*16+7],FIFO_12[256*6+x*16+7],FIFO_11[256*6+x*16+7],FIFO_10[256*6+x*16+7],FIFO_9[256*6+x*16+7],FIFO_8[256*6+x*16+7],FIFO_7[256*6+x*16+7],FIFO_6[256*6+x*16+7],FIFO_5[256*6+x*16+7],FIFO_4[256*6+x*16+7],FIFO_3[256*6+x*16+7],FIFO_2[256*6+x*16+7],FIFO_1[256*6+x*16+7],FIFO_16[256*7+x*16+7],FIFO_15[256*7+x*16+7],FIFO_14[256*7+x*16+7],FIFO_13[256*7+x*16+7],FIFO_12[256*7+x*16+7],FIFO_11[256*7+x*16+7],FIFO_10[256*7+x*16+7],FIFO_9[256*7+x*16+7],FIFO_8[256*7+x*16+7],FIFO_7[256*7+x*16+7],FIFO_6[256*7+x*16+7],FIFO_5[256*7+x*16+7],FIFO_4[256*7+x*16+7],FIFO_3[256*7+x*16+7],FIFO_2[256*7+x*16+7],FIFO_1[256*7+x*16+7],FIFO_16[256*8+x*16+7],FIFO_15[256*8+x*16+7],FIFO_14[256*8+x*16+7],FIFO_13[256*8+x*16+7],FIFO_12[256*8+x*16+7],FIFO_11[256*8+x*16+7],FIFO_10[256*8+x*16+7],FIFO_9[256*8+x*16+7],FIFO_8[256*8+x*16+7],FIFO_7[256*8+x*16+7],FIFO_6[256*8+x*16+7],FIFO_5[256*8+x*16+7],FIFO_4[256*8+x*16+7],FIFO_3[256*8+x*16+7],FIFO_2[256*8+x*16+7],FIFO_1[256*8+x*16+7],FIFO_16[256*9+x*16+7],FIFO_15[256*9+x*16+7],FIFO_14[256*9+x*16+7],FIFO_13[256*9+x*16+7],FIFO_12[256*9+x*16+7],FIFO_11[256*9+x*16+7],FIFO_10[256*9+x*16+7],FIFO_9[256*9+x*16+7],FIFO_8[256*9+x*16+7],FIFO_7[256*9+x*16+7],FIFO_6[256*9+x*16+7],FIFO_5[256*9+x*16+7],FIFO_4[256*9+x*16+7],FIFO_3[256*9+x*16+7],FIFO_2[256*9+x*16+7],FIFO_1[256*9+x*16+7],FIFO_16[256*10+x*16+7],FIFO_15[256*10+x*16+7],FIFO_14[256*10+x*16+7],FIFO_13[256*10+x*16+7],FIFO_12[256*10+x*16+7],FIFO_11[256*10+x*16+7],FIFO_10[256*10+x*16+7],FIFO_9[256*10+x*16+7],FIFO_8[256*10+x*16+7],FIFO_7[256*10+x*16+7],FIFO_6[256*10+x*16+7],FIFO_5[256*10+x*16+7],FIFO_4[256*10+x*16+7],FIFO_3[256*10+x*16+7],FIFO_2[256*10+x*16+7],FIFO_1[256*10+x*16+7],FIFO_16[256*11+x*16+7],FIFO_15[256*11+x*16+7],FIFO_14[256*11+x*16+7],FIFO_13[256*11+x*16+7],FIFO_12[256*11+x*16+7],FIFO_11[256*11+x*16+7],FIFO_10[256*11+x*16+7],FIFO_9[256*11+x*16+7],FIFO_8[256*11+x*16+7],FIFO_7[256*11+x*16+7],FIFO_6[256*11+x*16+7],FIFO_5[256*11+x*16+7],FIFO_4[256*11+x*16+7],FIFO_3[256*11+x*16+7],FIFO_2[256*11+x*16+7],FIFO_1[256*11+x*16+7],FIFO_16[256*12+x*16+7],FIFO_15[256*12+x*16+7],FIFO_14[256*12+x*16+7],FIFO_13[256*12+x*16+7],FIFO_12[256*12+x*16+7],FIFO_11[256*12+x*16+7],FIFO_10[256*12+x*16+7],FIFO_9[256*12+x*16+7],FIFO_8[256*12+x*16+7],FIFO_7[256*12+x*16+7],FIFO_6[256*12+x*16+7],FIFO_5[256*12+x*16+7],FIFO_4[256*12+x*16+7],FIFO_3[256*12+x*16+7],FIFO_2[256*12+x*16+7],FIFO_1[256*12+x*16+7],FIFO_16[256*13+x*16+7],FIFO_15[256*13+x*16+7],FIFO_14[256*13+x*16+7],FIFO_13[256*13+x*16+7],FIFO_12[256*13+x*16+7],FIFO_11[256*13+x*16+7],FIFO_10[256*13+x*16+7],FIFO_9[256*13+x*16+7],FIFO_8[256*13+x*16+7],FIFO_7[256*13+x*16+7],FIFO_6[256*13+x*16+7],FIFO_5[256*13+x*16+7],FIFO_4[256*13+x*16+7],FIFO_3[256*13+x*16+7],FIFO_2[256*13+x*16+7],FIFO_1[256*13+x*16+7],FIFO_16[256*14+x*16+7],FIFO_15[256*14+x*16+7],FIFO_14[256*14+x*16+7],FIFO_13[256*14+x*16+7],FIFO_12[256*14+x*16+7],FIFO_11[256*14+x*16+7],FIFO_10[256*14+x*16+7],FIFO_9[256*14+x*16+7],FIFO_8[256*14+x*16+7],FIFO_7[256*14+x*16+7],FIFO_6[256*14+x*16+7],FIFO_5[256*14+x*16+7],FIFO_4[256*14+x*16+7],FIFO_3[256*14+x*16+7],FIFO_2[256*14+x*16+7],FIFO_1[256*14+x*16+7],FIFO_16[256*15+x*16+7],FIFO_15[256*15+x*16+7],FIFO_14[256*15+x*16+7],FIFO_13[256*15+x*16+7],FIFO_12[256*15+x*16+7],FIFO_11[256*15+x*16+7],FIFO_10[256*15+x*16+7],FIFO_9[256*15+x*16+7],FIFO_8[256*15+x*16+7],FIFO_7[256*15+x*16+7],FIFO_6[256*15+x*16+7],FIFO_5[256*15+x*16+7],FIFO_4[256*15+x*16+7],FIFO_3[256*15+x*16+7],FIFO_2[256*15+x*16+7],FIFO_1[256*15+x*16+7]}; 
                error_vector9 <= dec9 ^ {FIFO_16[256*0+x*16+8],FIFO_15[256*0+x*16+8],FIFO_14[256*0+x*16+8],FIFO_13[256*0+x*16+8],FIFO_12[256*0+x*16+8],FIFO_11[256*0+x*16+8],FIFO_10[256*0+x*16+8],FIFO_9[256*0+x*16+8],FIFO_8[256*0+x*16+8],FIFO_7[256*0+x*16+8],FIFO_6[256*0+x*16+8],FIFO_5[256*0+x*16+8],FIFO_4[256*0+x*16+8],FIFO_3[256*0+x*16+8],FIFO_2[256*0+x*16+8],FIFO_1[256*0+x*16+8],FIFO_16[256*1+x*16+8],FIFO_15[256*1+x*16+8],FIFO_14[256*1+x*16+8],FIFO_13[256*1+x*16+8],FIFO_12[256*1+x*16+8],FIFO_11[256*1+x*16+8],FIFO_10[256*1+x*16+8],FIFO_9[256*1+x*16+8],FIFO_8[256*1+x*16+8],FIFO_7[256*1+x*16+8],FIFO_6[256*1+x*16+8],FIFO_5[256*1+x*16+8],FIFO_4[256*1+x*16+8],FIFO_3[256*1+x*16+8],FIFO_2[256*1+x*16+8],FIFO_1[256*1+x*16+8],FIFO_16[256*2+x*16+8],FIFO_15[256*2+x*16+8],FIFO_14[256*2+x*16+8],FIFO_13[256*2+x*16+8],FIFO_12[256*2+x*16+8],FIFO_11[256*2+x*16+8],FIFO_10[256*2+x*16+8],FIFO_9[256*2+x*16+8],FIFO_8[256*2+x*16+8],FIFO_7[256*2+x*16+8],FIFO_6[256*2+x*16+8],FIFO_5[256*2+x*16+8],FIFO_4[256*2+x*16+8],FIFO_3[256*2+x*16+8],FIFO_2[256*2+x*16+8],FIFO_1[256*2+x*16+8],FIFO_16[256*3+x*16+8],FIFO_15[256*3+x*16+8],FIFO_14[256*3+x*16+8],FIFO_13[256*3+x*16+8],FIFO_12[256*3+x*16+8],FIFO_11[256*3+x*16+8],FIFO_10[256*3+x*16+8],FIFO_9[256*3+x*16+8],FIFO_8[256*3+x*16+8],FIFO_7[256*3+x*16+8],FIFO_6[256*3+x*16+8],FIFO_5[256*3+x*16+8],FIFO_4[256*3+x*16+8],FIFO_3[256*3+x*16+8],FIFO_2[256*3+x*16+8],FIFO_1[256*3+x*16+8],FIFO_16[256*4+x*16+8],FIFO_15[256*4+x*16+8],FIFO_14[256*4+x*16+8],FIFO_13[256*4+x*16+8],FIFO_12[256*4+x*16+8],FIFO_11[256*4+x*16+8],FIFO_10[256*4+x*16+8],FIFO_9[256*4+x*16+8],FIFO_8[256*4+x*16+8],FIFO_7[256*4+x*16+8],FIFO_6[256*4+x*16+8],FIFO_5[256*4+x*16+8],FIFO_4[256*4+x*16+8],FIFO_3[256*4+x*16+8],FIFO_2[256*4+x*16+8],FIFO_1[256*4+x*16+8],FIFO_16[256*5+x*16+8],FIFO_15[256*5+x*16+8],FIFO_14[256*5+x*16+8],FIFO_13[256*5+x*16+8],FIFO_12[256*5+x*16+8],FIFO_11[256*5+x*16+8],FIFO_10[256*5+x*16+8],FIFO_9[256*5+x*16+8],FIFO_8[256*5+x*16+8],FIFO_7[256*5+x*16+8],FIFO_6[256*5+x*16+8],FIFO_5[256*5+x*16+8],FIFO_4[256*5+x*16+8],FIFO_3[256*5+x*16+8],FIFO_2[256*5+x*16+8],FIFO_1[256*5+x*16+8],FIFO_16[256*6+x*16+8],FIFO_15[256*6+x*16+8],FIFO_14[256*6+x*16+8],FIFO_13[256*6+x*16+8],FIFO_12[256*6+x*16+8],FIFO_11[256*6+x*16+8],FIFO_10[256*6+x*16+8],FIFO_9[256*6+x*16+8],FIFO_8[256*6+x*16+8],FIFO_7[256*6+x*16+8],FIFO_6[256*6+x*16+8],FIFO_5[256*6+x*16+8],FIFO_4[256*6+x*16+8],FIFO_3[256*6+x*16+8],FIFO_2[256*6+x*16+8],FIFO_1[256*6+x*16+8],FIFO_16[256*7+x*16+8],FIFO_15[256*7+x*16+8],FIFO_14[256*7+x*16+8],FIFO_13[256*7+x*16+8],FIFO_12[256*7+x*16+8],FIFO_11[256*7+x*16+8],FIFO_10[256*7+x*16+8],FIFO_9[256*7+x*16+8],FIFO_8[256*7+x*16+8],FIFO_7[256*7+x*16+8],FIFO_6[256*7+x*16+8],FIFO_5[256*7+x*16+8],FIFO_4[256*7+x*16+8],FIFO_3[256*7+x*16+8],FIFO_2[256*7+x*16+8],FIFO_1[256*7+x*16+8],FIFO_16[256*8+x*16+8],FIFO_15[256*8+x*16+8],FIFO_14[256*8+x*16+8],FIFO_13[256*8+x*16+8],FIFO_12[256*8+x*16+8],FIFO_11[256*8+x*16+8],FIFO_10[256*8+x*16+8],FIFO_9[256*8+x*16+8],FIFO_8[256*8+x*16+8],FIFO_7[256*8+x*16+8],FIFO_6[256*8+x*16+8],FIFO_5[256*8+x*16+8],FIFO_4[256*8+x*16+8],FIFO_3[256*8+x*16+8],FIFO_2[256*8+x*16+8],FIFO_1[256*8+x*16+8],FIFO_16[256*9+x*16+8],FIFO_15[256*9+x*16+8],FIFO_14[256*9+x*16+8],FIFO_13[256*9+x*16+8],FIFO_12[256*9+x*16+8],FIFO_11[256*9+x*16+8],FIFO_10[256*9+x*16+8],FIFO_9[256*9+x*16+8],FIFO_8[256*9+x*16+8],FIFO_7[256*9+x*16+8],FIFO_6[256*9+x*16+8],FIFO_5[256*9+x*16+8],FIFO_4[256*9+x*16+8],FIFO_3[256*9+x*16+8],FIFO_2[256*9+x*16+8],FIFO_1[256*9+x*16+8],FIFO_16[256*10+x*16+8],FIFO_15[256*10+x*16+8],FIFO_14[256*10+x*16+8],FIFO_13[256*10+x*16+8],FIFO_12[256*10+x*16+8],FIFO_11[256*10+x*16+8],FIFO_10[256*10+x*16+8],FIFO_9[256*10+x*16+8],FIFO_8[256*10+x*16+8],FIFO_7[256*10+x*16+8],FIFO_6[256*10+x*16+8],FIFO_5[256*10+x*16+8],FIFO_4[256*10+x*16+8],FIFO_3[256*10+x*16+8],FIFO_2[256*10+x*16+8],FIFO_1[256*10+x*16+8],FIFO_16[256*11+x*16+8],FIFO_15[256*11+x*16+8],FIFO_14[256*11+x*16+8],FIFO_13[256*11+x*16+8],FIFO_12[256*11+x*16+8],FIFO_11[256*11+x*16+8],FIFO_10[256*11+x*16+8],FIFO_9[256*11+x*16+8],FIFO_8[256*11+x*16+8],FIFO_7[256*11+x*16+8],FIFO_6[256*11+x*16+8],FIFO_5[256*11+x*16+8],FIFO_4[256*11+x*16+8],FIFO_3[256*11+x*16+8],FIFO_2[256*11+x*16+8],FIFO_1[256*11+x*16+8],FIFO_16[256*12+x*16+8],FIFO_15[256*12+x*16+8],FIFO_14[256*12+x*16+8],FIFO_13[256*12+x*16+8],FIFO_12[256*12+x*16+8],FIFO_11[256*12+x*16+8],FIFO_10[256*12+x*16+8],FIFO_9[256*12+x*16+8],FIFO_8[256*12+x*16+8],FIFO_7[256*12+x*16+8],FIFO_6[256*12+x*16+8],FIFO_5[256*12+x*16+8],FIFO_4[256*12+x*16+8],FIFO_3[256*12+x*16+8],FIFO_2[256*12+x*16+8],FIFO_1[256*12+x*16+8],FIFO_16[256*13+x*16+8],FIFO_15[256*13+x*16+8],FIFO_14[256*13+x*16+8],FIFO_13[256*13+x*16+8],FIFO_12[256*13+x*16+8],FIFO_11[256*13+x*16+8],FIFO_10[256*13+x*16+8],FIFO_9[256*13+x*16+8],FIFO_8[256*13+x*16+8],FIFO_7[256*13+x*16+8],FIFO_6[256*13+x*16+8],FIFO_5[256*13+x*16+8],FIFO_4[256*13+x*16+8],FIFO_3[256*13+x*16+8],FIFO_2[256*13+x*16+8],FIFO_1[256*13+x*16+8],FIFO_16[256*14+x*16+8],FIFO_15[256*14+x*16+8],FIFO_14[256*14+x*16+8],FIFO_13[256*14+x*16+8],FIFO_12[256*14+x*16+8],FIFO_11[256*14+x*16+8],FIFO_10[256*14+x*16+8],FIFO_9[256*14+x*16+8],FIFO_8[256*14+x*16+8],FIFO_7[256*14+x*16+8],FIFO_6[256*14+x*16+8],FIFO_5[256*14+x*16+8],FIFO_4[256*14+x*16+8],FIFO_3[256*14+x*16+8],FIFO_2[256*14+x*16+8],FIFO_1[256*14+x*16+8],FIFO_16[256*15+x*16+8],FIFO_15[256*15+x*16+8],FIFO_14[256*15+x*16+8],FIFO_13[256*15+x*16+8],FIFO_12[256*15+x*16+8],FIFO_11[256*15+x*16+8],FIFO_10[256*15+x*16+8],FIFO_9[256*15+x*16+8],FIFO_8[256*15+x*16+8],FIFO_7[256*15+x*16+8],FIFO_6[256*15+x*16+8],FIFO_5[256*15+x*16+8],FIFO_4[256*15+x*16+8],FIFO_3[256*15+x*16+8],FIFO_2[256*15+x*16+8],FIFO_1[256*15+x*16+8]}; 
                error_vector10 <= dec10 ^ {FIFO_16[256*0+x*16+9],FIFO_15[256*0+x*16+9],FIFO_14[256*0+x*16+9],FIFO_13[256*0+x*16+9],FIFO_12[256*0+x*16+9],FIFO_11[256*0+x*16+9],FIFO_10[256*0+x*16+9],FIFO_9[256*0+x*16+9],FIFO_8[256*0+x*16+9],FIFO_7[256*0+x*16+9],FIFO_6[256*0+x*16+9],FIFO_5[256*0+x*16+9],FIFO_4[256*0+x*16+9],FIFO_3[256*0+x*16+9],FIFO_2[256*0+x*16+9],FIFO_1[256*0+x*16+9],FIFO_16[256*1+x*16+9],FIFO_15[256*1+x*16+9],FIFO_14[256*1+x*16+9],FIFO_13[256*1+x*16+9],FIFO_12[256*1+x*16+9],FIFO_11[256*1+x*16+9],FIFO_10[256*1+x*16+9],FIFO_9[256*1+x*16+9],FIFO_8[256*1+x*16+9],FIFO_7[256*1+x*16+9],FIFO_6[256*1+x*16+9],FIFO_5[256*1+x*16+9],FIFO_4[256*1+x*16+9],FIFO_3[256*1+x*16+9],FIFO_2[256*1+x*16+9],FIFO_1[256*1+x*16+9],FIFO_16[256*2+x*16+9],FIFO_15[256*2+x*16+9],FIFO_14[256*2+x*16+9],FIFO_13[256*2+x*16+9],FIFO_12[256*2+x*16+9],FIFO_11[256*2+x*16+9],FIFO_10[256*2+x*16+9],FIFO_9[256*2+x*16+9],FIFO_8[256*2+x*16+9],FIFO_7[256*2+x*16+9],FIFO_6[256*2+x*16+9],FIFO_5[256*2+x*16+9],FIFO_4[256*2+x*16+9],FIFO_3[256*2+x*16+9],FIFO_2[256*2+x*16+9],FIFO_1[256*2+x*16+9],FIFO_16[256*3+x*16+9],FIFO_15[256*3+x*16+9],FIFO_14[256*3+x*16+9],FIFO_13[256*3+x*16+9],FIFO_12[256*3+x*16+9],FIFO_11[256*3+x*16+9],FIFO_10[256*3+x*16+9],FIFO_9[256*3+x*16+9],FIFO_8[256*3+x*16+9],FIFO_7[256*3+x*16+9],FIFO_6[256*3+x*16+9],FIFO_5[256*3+x*16+9],FIFO_4[256*3+x*16+9],FIFO_3[256*3+x*16+9],FIFO_2[256*3+x*16+9],FIFO_1[256*3+x*16+9],FIFO_16[256*4+x*16+9],FIFO_15[256*4+x*16+9],FIFO_14[256*4+x*16+9],FIFO_13[256*4+x*16+9],FIFO_12[256*4+x*16+9],FIFO_11[256*4+x*16+9],FIFO_10[256*4+x*16+9],FIFO_9[256*4+x*16+9],FIFO_8[256*4+x*16+9],FIFO_7[256*4+x*16+9],FIFO_6[256*4+x*16+9],FIFO_5[256*4+x*16+9],FIFO_4[256*4+x*16+9],FIFO_3[256*4+x*16+9],FIFO_2[256*4+x*16+9],FIFO_1[256*4+x*16+9],FIFO_16[256*5+x*16+9],FIFO_15[256*5+x*16+9],FIFO_14[256*5+x*16+9],FIFO_13[256*5+x*16+9],FIFO_12[256*5+x*16+9],FIFO_11[256*5+x*16+9],FIFO_10[256*5+x*16+9],FIFO_9[256*5+x*16+9],FIFO_8[256*5+x*16+9],FIFO_7[256*5+x*16+9],FIFO_6[256*5+x*16+9],FIFO_5[256*5+x*16+9],FIFO_4[256*5+x*16+9],FIFO_3[256*5+x*16+9],FIFO_2[256*5+x*16+9],FIFO_1[256*5+x*16+9],FIFO_16[256*6+x*16+9],FIFO_15[256*6+x*16+9],FIFO_14[256*6+x*16+9],FIFO_13[256*6+x*16+9],FIFO_12[256*6+x*16+9],FIFO_11[256*6+x*16+9],FIFO_10[256*6+x*16+9],FIFO_9[256*6+x*16+9],FIFO_8[256*6+x*16+9],FIFO_7[256*6+x*16+9],FIFO_6[256*6+x*16+9],FIFO_5[256*6+x*16+9],FIFO_4[256*6+x*16+9],FIFO_3[256*6+x*16+9],FIFO_2[256*6+x*16+9],FIFO_1[256*6+x*16+9],FIFO_16[256*7+x*16+9],FIFO_15[256*7+x*16+9],FIFO_14[256*7+x*16+9],FIFO_13[256*7+x*16+9],FIFO_12[256*7+x*16+9],FIFO_11[256*7+x*16+9],FIFO_10[256*7+x*16+9],FIFO_9[256*7+x*16+9],FIFO_8[256*7+x*16+9],FIFO_7[256*7+x*16+9],FIFO_6[256*7+x*16+9],FIFO_5[256*7+x*16+9],FIFO_4[256*7+x*16+9],FIFO_3[256*7+x*16+9],FIFO_2[256*7+x*16+9],FIFO_1[256*7+x*16+9],FIFO_16[256*8+x*16+9],FIFO_15[256*8+x*16+9],FIFO_14[256*8+x*16+9],FIFO_13[256*8+x*16+9],FIFO_12[256*8+x*16+9],FIFO_11[256*8+x*16+9],FIFO_10[256*8+x*16+9],FIFO_9[256*8+x*16+9],FIFO_8[256*8+x*16+9],FIFO_7[256*8+x*16+9],FIFO_6[256*8+x*16+9],FIFO_5[256*8+x*16+9],FIFO_4[256*8+x*16+9],FIFO_3[256*8+x*16+9],FIFO_2[256*8+x*16+9],FIFO_1[256*8+x*16+9],FIFO_16[256*9+x*16+9],FIFO_15[256*9+x*16+9],FIFO_14[256*9+x*16+9],FIFO_13[256*9+x*16+9],FIFO_12[256*9+x*16+9],FIFO_11[256*9+x*16+9],FIFO_10[256*9+x*16+9],FIFO_9[256*9+x*16+9],FIFO_8[256*9+x*16+9],FIFO_7[256*9+x*16+9],FIFO_6[256*9+x*16+9],FIFO_5[256*9+x*16+9],FIFO_4[256*9+x*16+9],FIFO_3[256*9+x*16+9],FIFO_2[256*9+x*16+9],FIFO_1[256*9+x*16+9],FIFO_16[256*10+x*16+9],FIFO_15[256*10+x*16+9],FIFO_14[256*10+x*16+9],FIFO_13[256*10+x*16+9],FIFO_12[256*10+x*16+9],FIFO_11[256*10+x*16+9],FIFO_10[256*10+x*16+9],FIFO_9[256*10+x*16+9],FIFO_8[256*10+x*16+9],FIFO_7[256*10+x*16+9],FIFO_6[256*10+x*16+9],FIFO_5[256*10+x*16+9],FIFO_4[256*10+x*16+9],FIFO_3[256*10+x*16+9],FIFO_2[256*10+x*16+9],FIFO_1[256*10+x*16+9],FIFO_16[256*11+x*16+9],FIFO_15[256*11+x*16+9],FIFO_14[256*11+x*16+9],FIFO_13[256*11+x*16+9],FIFO_12[256*11+x*16+9],FIFO_11[256*11+x*16+9],FIFO_10[256*11+x*16+9],FIFO_9[256*11+x*16+9],FIFO_8[256*11+x*16+9],FIFO_7[256*11+x*16+9],FIFO_6[256*11+x*16+9],FIFO_5[256*11+x*16+9],FIFO_4[256*11+x*16+9],FIFO_3[256*11+x*16+9],FIFO_2[256*11+x*16+9],FIFO_1[256*11+x*16+9],FIFO_16[256*12+x*16+9],FIFO_15[256*12+x*16+9],FIFO_14[256*12+x*16+9],FIFO_13[256*12+x*16+9],FIFO_12[256*12+x*16+9],FIFO_11[256*12+x*16+9],FIFO_10[256*12+x*16+9],FIFO_9[256*12+x*16+9],FIFO_8[256*12+x*16+9],FIFO_7[256*12+x*16+9],FIFO_6[256*12+x*16+9],FIFO_5[256*12+x*16+9],FIFO_4[256*12+x*16+9],FIFO_3[256*12+x*16+9],FIFO_2[256*12+x*16+9],FIFO_1[256*12+x*16+9],FIFO_16[256*13+x*16+9],FIFO_15[256*13+x*16+9],FIFO_14[256*13+x*16+9],FIFO_13[256*13+x*16+9],FIFO_12[256*13+x*16+9],FIFO_11[256*13+x*16+9],FIFO_10[256*13+x*16+9],FIFO_9[256*13+x*16+9],FIFO_8[256*13+x*16+9],FIFO_7[256*13+x*16+9],FIFO_6[256*13+x*16+9],FIFO_5[256*13+x*16+9],FIFO_4[256*13+x*16+9],FIFO_3[256*13+x*16+9],FIFO_2[256*13+x*16+9],FIFO_1[256*13+x*16+9],FIFO_16[256*14+x*16+9],FIFO_15[256*14+x*16+9],FIFO_14[256*14+x*16+9],FIFO_13[256*14+x*16+9],FIFO_12[256*14+x*16+9],FIFO_11[256*14+x*16+9],FIFO_10[256*14+x*16+9],FIFO_9[256*14+x*16+9],FIFO_8[256*14+x*16+9],FIFO_7[256*14+x*16+9],FIFO_6[256*14+x*16+9],FIFO_5[256*14+x*16+9],FIFO_4[256*14+x*16+9],FIFO_3[256*14+x*16+9],FIFO_2[256*14+x*16+9],FIFO_1[256*14+x*16+9],FIFO_16[256*15+x*16+9],FIFO_15[256*15+x*16+9],FIFO_14[256*15+x*16+9],FIFO_13[256*15+x*16+9],FIFO_12[256*15+x*16+9],FIFO_11[256*15+x*16+9],FIFO_10[256*15+x*16+9],FIFO_9[256*15+x*16+9],FIFO_8[256*15+x*16+9],FIFO_7[256*15+x*16+9],FIFO_6[256*15+x*16+9],FIFO_5[256*15+x*16+9],FIFO_4[256*15+x*16+9],FIFO_3[256*15+x*16+9],FIFO_2[256*15+x*16+9],FIFO_1[256*15+x*16+9]}; 
                error_vector11 <= dec11 ^ {FIFO_16[256*0+x*16+10],FIFO_15[256*0+x*16+10],FIFO_14[256*0+x*16+10],FIFO_13[256*0+x*16+10],FIFO_12[256*0+x*16+10],FIFO_11[256*0+x*16+10],FIFO_10[256*0+x*16+10],FIFO_9[256*0+x*16+10],FIFO_8[256*0+x*16+10],FIFO_7[256*0+x*16+10],FIFO_6[256*0+x*16+10],FIFO_5[256*0+x*16+10],FIFO_4[256*0+x*16+10],FIFO_3[256*0+x*16+10],FIFO_2[256*0+x*16+10],FIFO_1[256*0+x*16+10],FIFO_16[256*1+x*16+10],FIFO_15[256*1+x*16+10],FIFO_14[256*1+x*16+10],FIFO_13[256*1+x*16+10],FIFO_12[256*1+x*16+10],FIFO_11[256*1+x*16+10],FIFO_10[256*1+x*16+10],FIFO_9[256*1+x*16+10],FIFO_8[256*1+x*16+10],FIFO_7[256*1+x*16+10],FIFO_6[256*1+x*16+10],FIFO_5[256*1+x*16+10],FIFO_4[256*1+x*16+10],FIFO_3[256*1+x*16+10],FIFO_2[256*1+x*16+10],FIFO_1[256*1+x*16+10],FIFO_16[256*2+x*16+10],FIFO_15[256*2+x*16+10],FIFO_14[256*2+x*16+10],FIFO_13[256*2+x*16+10],FIFO_12[256*2+x*16+10],FIFO_11[256*2+x*16+10],FIFO_10[256*2+x*16+10],FIFO_9[256*2+x*16+10],FIFO_8[256*2+x*16+10],FIFO_7[256*2+x*16+10],FIFO_6[256*2+x*16+10],FIFO_5[256*2+x*16+10],FIFO_4[256*2+x*16+10],FIFO_3[256*2+x*16+10],FIFO_2[256*2+x*16+10],FIFO_1[256*2+x*16+10],FIFO_16[256*3+x*16+10],FIFO_15[256*3+x*16+10],FIFO_14[256*3+x*16+10],FIFO_13[256*3+x*16+10],FIFO_12[256*3+x*16+10],FIFO_11[256*3+x*16+10],FIFO_10[256*3+x*16+10],FIFO_9[256*3+x*16+10],FIFO_8[256*3+x*16+10],FIFO_7[256*3+x*16+10],FIFO_6[256*3+x*16+10],FIFO_5[256*3+x*16+10],FIFO_4[256*3+x*16+10],FIFO_3[256*3+x*16+10],FIFO_2[256*3+x*16+10],FIFO_1[256*3+x*16+10],FIFO_16[256*4+x*16+10],FIFO_15[256*4+x*16+10],FIFO_14[256*4+x*16+10],FIFO_13[256*4+x*16+10],FIFO_12[256*4+x*16+10],FIFO_11[256*4+x*16+10],FIFO_10[256*4+x*16+10],FIFO_9[256*4+x*16+10],FIFO_8[256*4+x*16+10],FIFO_7[256*4+x*16+10],FIFO_6[256*4+x*16+10],FIFO_5[256*4+x*16+10],FIFO_4[256*4+x*16+10],FIFO_3[256*4+x*16+10],FIFO_2[256*4+x*16+10],FIFO_1[256*4+x*16+10],FIFO_16[256*5+x*16+10],FIFO_15[256*5+x*16+10],FIFO_14[256*5+x*16+10],FIFO_13[256*5+x*16+10],FIFO_12[256*5+x*16+10],FIFO_11[256*5+x*16+10],FIFO_10[256*5+x*16+10],FIFO_9[256*5+x*16+10],FIFO_8[256*5+x*16+10],FIFO_7[256*5+x*16+10],FIFO_6[256*5+x*16+10],FIFO_5[256*5+x*16+10],FIFO_4[256*5+x*16+10],FIFO_3[256*5+x*16+10],FIFO_2[256*5+x*16+10],FIFO_1[256*5+x*16+10],FIFO_16[256*6+x*16+10],FIFO_15[256*6+x*16+10],FIFO_14[256*6+x*16+10],FIFO_13[256*6+x*16+10],FIFO_12[256*6+x*16+10],FIFO_11[256*6+x*16+10],FIFO_10[256*6+x*16+10],FIFO_9[256*6+x*16+10],FIFO_8[256*6+x*16+10],FIFO_7[256*6+x*16+10],FIFO_6[256*6+x*16+10],FIFO_5[256*6+x*16+10],FIFO_4[256*6+x*16+10],FIFO_3[256*6+x*16+10],FIFO_2[256*6+x*16+10],FIFO_1[256*6+x*16+10],FIFO_16[256*7+x*16+10],FIFO_15[256*7+x*16+10],FIFO_14[256*7+x*16+10],FIFO_13[256*7+x*16+10],FIFO_12[256*7+x*16+10],FIFO_11[256*7+x*16+10],FIFO_10[256*7+x*16+10],FIFO_9[256*7+x*16+10],FIFO_8[256*7+x*16+10],FIFO_7[256*7+x*16+10],FIFO_6[256*7+x*16+10],FIFO_5[256*7+x*16+10],FIFO_4[256*7+x*16+10],FIFO_3[256*7+x*16+10],FIFO_2[256*7+x*16+10],FIFO_1[256*7+x*16+10],FIFO_16[256*8+x*16+10],FIFO_15[256*8+x*16+10],FIFO_14[256*8+x*16+10],FIFO_13[256*8+x*16+10],FIFO_12[256*8+x*16+10],FIFO_11[256*8+x*16+10],FIFO_10[256*8+x*16+10],FIFO_9[256*8+x*16+10],FIFO_8[256*8+x*16+10],FIFO_7[256*8+x*16+10],FIFO_6[256*8+x*16+10],FIFO_5[256*8+x*16+10],FIFO_4[256*8+x*16+10],FIFO_3[256*8+x*16+10],FIFO_2[256*8+x*16+10],FIFO_1[256*8+x*16+10],FIFO_16[256*9+x*16+10],FIFO_15[256*9+x*16+10],FIFO_14[256*9+x*16+10],FIFO_13[256*9+x*16+10],FIFO_12[256*9+x*16+10],FIFO_11[256*9+x*16+10],FIFO_10[256*9+x*16+10],FIFO_9[256*9+x*16+10],FIFO_8[256*9+x*16+10],FIFO_7[256*9+x*16+10],FIFO_6[256*9+x*16+10],FIFO_5[256*9+x*16+10],FIFO_4[256*9+x*16+10],FIFO_3[256*9+x*16+10],FIFO_2[256*9+x*16+10],FIFO_1[256*9+x*16+10],FIFO_16[256*10+x*16+10],FIFO_15[256*10+x*16+10],FIFO_14[256*10+x*16+10],FIFO_13[256*10+x*16+10],FIFO_12[256*10+x*16+10],FIFO_11[256*10+x*16+10],FIFO_10[256*10+x*16+10],FIFO_9[256*10+x*16+10],FIFO_8[256*10+x*16+10],FIFO_7[256*10+x*16+10],FIFO_6[256*10+x*16+10],FIFO_5[256*10+x*16+10],FIFO_4[256*10+x*16+10],FIFO_3[256*10+x*16+10],FIFO_2[256*10+x*16+10],FIFO_1[256*10+x*16+10],FIFO_16[256*11+x*16+10],FIFO_15[256*11+x*16+10],FIFO_14[256*11+x*16+10],FIFO_13[256*11+x*16+10],FIFO_12[256*11+x*16+10],FIFO_11[256*11+x*16+10],FIFO_10[256*11+x*16+10],FIFO_9[256*11+x*16+10],FIFO_8[256*11+x*16+10],FIFO_7[256*11+x*16+10],FIFO_6[256*11+x*16+10],FIFO_5[256*11+x*16+10],FIFO_4[256*11+x*16+10],FIFO_3[256*11+x*16+10],FIFO_2[256*11+x*16+10],FIFO_1[256*11+x*16+10],FIFO_16[256*12+x*16+10],FIFO_15[256*12+x*16+10],FIFO_14[256*12+x*16+10],FIFO_13[256*12+x*16+10],FIFO_12[256*12+x*16+10],FIFO_11[256*12+x*16+10],FIFO_10[256*12+x*16+10],FIFO_9[256*12+x*16+10],FIFO_8[256*12+x*16+10],FIFO_7[256*12+x*16+10],FIFO_6[256*12+x*16+10],FIFO_5[256*12+x*16+10],FIFO_4[256*12+x*16+10],FIFO_3[256*12+x*16+10],FIFO_2[256*12+x*16+10],FIFO_1[256*12+x*16+10],FIFO_16[256*13+x*16+10],FIFO_15[256*13+x*16+10],FIFO_14[256*13+x*16+10],FIFO_13[256*13+x*16+10],FIFO_12[256*13+x*16+10],FIFO_11[256*13+x*16+10],FIFO_10[256*13+x*16+10],FIFO_9[256*13+x*16+10],FIFO_8[256*13+x*16+10],FIFO_7[256*13+x*16+10],FIFO_6[256*13+x*16+10],FIFO_5[256*13+x*16+10],FIFO_4[256*13+x*16+10],FIFO_3[256*13+x*16+10],FIFO_2[256*13+x*16+10],FIFO_1[256*13+x*16+10],FIFO_16[256*14+x*16+10],FIFO_15[256*14+x*16+10],FIFO_14[256*14+x*16+10],FIFO_13[256*14+x*16+10],FIFO_12[256*14+x*16+10],FIFO_11[256*14+x*16+10],FIFO_10[256*14+x*16+10],FIFO_9[256*14+x*16+10],FIFO_8[256*14+x*16+10],FIFO_7[256*14+x*16+10],FIFO_6[256*14+x*16+10],FIFO_5[256*14+x*16+10],FIFO_4[256*14+x*16+10],FIFO_3[256*14+x*16+10],FIFO_2[256*14+x*16+10],FIFO_1[256*14+x*16+10],FIFO_16[256*15+x*16+10],FIFO_15[256*15+x*16+10],FIFO_14[256*15+x*16+10],FIFO_13[256*15+x*16+10],FIFO_12[256*15+x*16+10],FIFO_11[256*15+x*16+10],FIFO_10[256*15+x*16+10],FIFO_9[256*15+x*16+10],FIFO_8[256*15+x*16+10],FIFO_7[256*15+x*16+10],FIFO_6[256*15+x*16+10],FIFO_5[256*15+x*16+10],FIFO_4[256*15+x*16+10],FIFO_3[256*15+x*16+10],FIFO_2[256*15+x*16+10],FIFO_1[256*15+x*16+10]}; 
                error_vector12 <= dec12 ^ {FIFO_16[256*0+x*16+11],FIFO_15[256*0+x*16+11],FIFO_14[256*0+x*16+11],FIFO_13[256*0+x*16+11],FIFO_12[256*0+x*16+11],FIFO_11[256*0+x*16+11],FIFO_10[256*0+x*16+11],FIFO_9[256*0+x*16+11],FIFO_8[256*0+x*16+11],FIFO_7[256*0+x*16+11],FIFO_6[256*0+x*16+11],FIFO_5[256*0+x*16+11],FIFO_4[256*0+x*16+11],FIFO_3[256*0+x*16+11],FIFO_2[256*0+x*16+11],FIFO_1[256*0+x*16+11],FIFO_16[256*1+x*16+11],FIFO_15[256*1+x*16+11],FIFO_14[256*1+x*16+11],FIFO_13[256*1+x*16+11],FIFO_12[256*1+x*16+11],FIFO_11[256*1+x*16+11],FIFO_10[256*1+x*16+11],FIFO_9[256*1+x*16+11],FIFO_8[256*1+x*16+11],FIFO_7[256*1+x*16+11],FIFO_6[256*1+x*16+11],FIFO_5[256*1+x*16+11],FIFO_4[256*1+x*16+11],FIFO_3[256*1+x*16+11],FIFO_2[256*1+x*16+11],FIFO_1[256*1+x*16+11],FIFO_16[256*2+x*16+11],FIFO_15[256*2+x*16+11],FIFO_14[256*2+x*16+11],FIFO_13[256*2+x*16+11],FIFO_12[256*2+x*16+11],FIFO_11[256*2+x*16+11],FIFO_10[256*2+x*16+11],FIFO_9[256*2+x*16+11],FIFO_8[256*2+x*16+11],FIFO_7[256*2+x*16+11],FIFO_6[256*2+x*16+11],FIFO_5[256*2+x*16+11],FIFO_4[256*2+x*16+11],FIFO_3[256*2+x*16+11],FIFO_2[256*2+x*16+11],FIFO_1[256*2+x*16+11],FIFO_16[256*3+x*16+11],FIFO_15[256*3+x*16+11],FIFO_14[256*3+x*16+11],FIFO_13[256*3+x*16+11],FIFO_12[256*3+x*16+11],FIFO_11[256*3+x*16+11],FIFO_10[256*3+x*16+11],FIFO_9[256*3+x*16+11],FIFO_8[256*3+x*16+11],FIFO_7[256*3+x*16+11],FIFO_6[256*3+x*16+11],FIFO_5[256*3+x*16+11],FIFO_4[256*3+x*16+11],FIFO_3[256*3+x*16+11],FIFO_2[256*3+x*16+11],FIFO_1[256*3+x*16+11],FIFO_16[256*4+x*16+11],FIFO_15[256*4+x*16+11],FIFO_14[256*4+x*16+11],FIFO_13[256*4+x*16+11],FIFO_12[256*4+x*16+11],FIFO_11[256*4+x*16+11],FIFO_10[256*4+x*16+11],FIFO_9[256*4+x*16+11],FIFO_8[256*4+x*16+11],FIFO_7[256*4+x*16+11],FIFO_6[256*4+x*16+11],FIFO_5[256*4+x*16+11],FIFO_4[256*4+x*16+11],FIFO_3[256*4+x*16+11],FIFO_2[256*4+x*16+11],FIFO_1[256*4+x*16+11],FIFO_16[256*5+x*16+11],FIFO_15[256*5+x*16+11],FIFO_14[256*5+x*16+11],FIFO_13[256*5+x*16+11],FIFO_12[256*5+x*16+11],FIFO_11[256*5+x*16+11],FIFO_10[256*5+x*16+11],FIFO_9[256*5+x*16+11],FIFO_8[256*5+x*16+11],FIFO_7[256*5+x*16+11],FIFO_6[256*5+x*16+11],FIFO_5[256*5+x*16+11],FIFO_4[256*5+x*16+11],FIFO_3[256*5+x*16+11],FIFO_2[256*5+x*16+11],FIFO_1[256*5+x*16+11],FIFO_16[256*6+x*16+11],FIFO_15[256*6+x*16+11],FIFO_14[256*6+x*16+11],FIFO_13[256*6+x*16+11],FIFO_12[256*6+x*16+11],FIFO_11[256*6+x*16+11],FIFO_10[256*6+x*16+11],FIFO_9[256*6+x*16+11],FIFO_8[256*6+x*16+11],FIFO_7[256*6+x*16+11],FIFO_6[256*6+x*16+11],FIFO_5[256*6+x*16+11],FIFO_4[256*6+x*16+11],FIFO_3[256*6+x*16+11],FIFO_2[256*6+x*16+11],FIFO_1[256*6+x*16+11],FIFO_16[256*7+x*16+11],FIFO_15[256*7+x*16+11],FIFO_14[256*7+x*16+11],FIFO_13[256*7+x*16+11],FIFO_12[256*7+x*16+11],FIFO_11[256*7+x*16+11],FIFO_10[256*7+x*16+11],FIFO_9[256*7+x*16+11],FIFO_8[256*7+x*16+11],FIFO_7[256*7+x*16+11],FIFO_6[256*7+x*16+11],FIFO_5[256*7+x*16+11],FIFO_4[256*7+x*16+11],FIFO_3[256*7+x*16+11],FIFO_2[256*7+x*16+11],FIFO_1[256*7+x*16+11],FIFO_16[256*8+x*16+11],FIFO_15[256*8+x*16+11],FIFO_14[256*8+x*16+11],FIFO_13[256*8+x*16+11],FIFO_12[256*8+x*16+11],FIFO_11[256*8+x*16+11],FIFO_10[256*8+x*16+11],FIFO_9[256*8+x*16+11],FIFO_8[256*8+x*16+11],FIFO_7[256*8+x*16+11],FIFO_6[256*8+x*16+11],FIFO_5[256*8+x*16+11],FIFO_4[256*8+x*16+11],FIFO_3[256*8+x*16+11],FIFO_2[256*8+x*16+11],FIFO_1[256*8+x*16+11],FIFO_16[256*9+x*16+11],FIFO_15[256*9+x*16+11],FIFO_14[256*9+x*16+11],FIFO_13[256*9+x*16+11],FIFO_12[256*9+x*16+11],FIFO_11[256*9+x*16+11],FIFO_10[256*9+x*16+11],FIFO_9[256*9+x*16+11],FIFO_8[256*9+x*16+11],FIFO_7[256*9+x*16+11],FIFO_6[256*9+x*16+11],FIFO_5[256*9+x*16+11],FIFO_4[256*9+x*16+11],FIFO_3[256*9+x*16+11],FIFO_2[256*9+x*16+11],FIFO_1[256*9+x*16+11],FIFO_16[256*10+x*16+11],FIFO_15[256*10+x*16+11],FIFO_14[256*10+x*16+11],FIFO_13[256*10+x*16+11],FIFO_12[256*10+x*16+11],FIFO_11[256*10+x*16+11],FIFO_10[256*10+x*16+11],FIFO_9[256*10+x*16+11],FIFO_8[256*10+x*16+11],FIFO_7[256*10+x*16+11],FIFO_6[256*10+x*16+11],FIFO_5[256*10+x*16+11],FIFO_4[256*10+x*16+11],FIFO_3[256*10+x*16+11],FIFO_2[256*10+x*16+11],FIFO_1[256*10+x*16+11],FIFO_16[256*11+x*16+11],FIFO_15[256*11+x*16+11],FIFO_14[256*11+x*16+11],FIFO_13[256*11+x*16+11],FIFO_12[256*11+x*16+11],FIFO_11[256*11+x*16+11],FIFO_10[256*11+x*16+11],FIFO_9[256*11+x*16+11],FIFO_8[256*11+x*16+11],FIFO_7[256*11+x*16+11],FIFO_6[256*11+x*16+11],FIFO_5[256*11+x*16+11],FIFO_4[256*11+x*16+11],FIFO_3[256*11+x*16+11],FIFO_2[256*11+x*16+11],FIFO_1[256*11+x*16+11],FIFO_16[256*12+x*16+11],FIFO_15[256*12+x*16+11],FIFO_14[256*12+x*16+11],FIFO_13[256*12+x*16+11],FIFO_12[256*12+x*16+11],FIFO_11[256*12+x*16+11],FIFO_10[256*12+x*16+11],FIFO_9[256*12+x*16+11],FIFO_8[256*12+x*16+11],FIFO_7[256*12+x*16+11],FIFO_6[256*12+x*16+11],FIFO_5[256*12+x*16+11],FIFO_4[256*12+x*16+11],FIFO_3[256*12+x*16+11],FIFO_2[256*12+x*16+11],FIFO_1[256*12+x*16+11],FIFO_16[256*13+x*16+11],FIFO_15[256*13+x*16+11],FIFO_14[256*13+x*16+11],FIFO_13[256*13+x*16+11],FIFO_12[256*13+x*16+11],FIFO_11[256*13+x*16+11],FIFO_10[256*13+x*16+11],FIFO_9[256*13+x*16+11],FIFO_8[256*13+x*16+11],FIFO_7[256*13+x*16+11],FIFO_6[256*13+x*16+11],FIFO_5[256*13+x*16+11],FIFO_4[256*13+x*16+11],FIFO_3[256*13+x*16+11],FIFO_2[256*13+x*16+11],FIFO_1[256*13+x*16+11],FIFO_16[256*14+x*16+11],FIFO_15[256*14+x*16+11],FIFO_14[256*14+x*16+11],FIFO_13[256*14+x*16+11],FIFO_12[256*14+x*16+11],FIFO_11[256*14+x*16+11],FIFO_10[256*14+x*16+11],FIFO_9[256*14+x*16+11],FIFO_8[256*14+x*16+11],FIFO_7[256*14+x*16+11],FIFO_6[256*14+x*16+11],FIFO_5[256*14+x*16+11],FIFO_4[256*14+x*16+11],FIFO_3[256*14+x*16+11],FIFO_2[256*14+x*16+11],FIFO_1[256*14+x*16+11],FIFO_16[256*15+x*16+11],FIFO_15[256*15+x*16+11],FIFO_14[256*15+x*16+11],FIFO_13[256*15+x*16+11],FIFO_12[256*15+x*16+11],FIFO_11[256*15+x*16+11],FIFO_10[256*15+x*16+11],FIFO_9[256*15+x*16+11],FIFO_8[256*15+x*16+11],FIFO_7[256*15+x*16+11],FIFO_6[256*15+x*16+11],FIFO_5[256*15+x*16+11],FIFO_4[256*15+x*16+11],FIFO_3[256*15+x*16+11],FIFO_2[256*15+x*16+11],FIFO_1[256*15+x*16+11]}; 
                error_vector13 <= dec13 ^ {FIFO_16[256*0+x*16+12],FIFO_15[256*0+x*16+12],FIFO_14[256*0+x*16+12],FIFO_13[256*0+x*16+12],FIFO_12[256*0+x*16+12],FIFO_11[256*0+x*16+12],FIFO_10[256*0+x*16+12],FIFO_9[256*0+x*16+12],FIFO_8[256*0+x*16+12],FIFO_7[256*0+x*16+12],FIFO_6[256*0+x*16+12],FIFO_5[256*0+x*16+12],FIFO_4[256*0+x*16+12],FIFO_3[256*0+x*16+12],FIFO_2[256*0+x*16+12],FIFO_1[256*0+x*16+12],FIFO_16[256*1+x*16+12],FIFO_15[256*1+x*16+12],FIFO_14[256*1+x*16+12],FIFO_13[256*1+x*16+12],FIFO_12[256*1+x*16+12],FIFO_11[256*1+x*16+12],FIFO_10[256*1+x*16+12],FIFO_9[256*1+x*16+12],FIFO_8[256*1+x*16+12],FIFO_7[256*1+x*16+12],FIFO_6[256*1+x*16+12],FIFO_5[256*1+x*16+12],FIFO_4[256*1+x*16+12],FIFO_3[256*1+x*16+12],FIFO_2[256*1+x*16+12],FIFO_1[256*1+x*16+12],FIFO_16[256*2+x*16+12],FIFO_15[256*2+x*16+12],FIFO_14[256*2+x*16+12],FIFO_13[256*2+x*16+12],FIFO_12[256*2+x*16+12],FIFO_11[256*2+x*16+12],FIFO_10[256*2+x*16+12],FIFO_9[256*2+x*16+12],FIFO_8[256*2+x*16+12],FIFO_7[256*2+x*16+12],FIFO_6[256*2+x*16+12],FIFO_5[256*2+x*16+12],FIFO_4[256*2+x*16+12],FIFO_3[256*2+x*16+12],FIFO_2[256*2+x*16+12],FIFO_1[256*2+x*16+12],FIFO_16[256*3+x*16+12],FIFO_15[256*3+x*16+12],FIFO_14[256*3+x*16+12],FIFO_13[256*3+x*16+12],FIFO_12[256*3+x*16+12],FIFO_11[256*3+x*16+12],FIFO_10[256*3+x*16+12],FIFO_9[256*3+x*16+12],FIFO_8[256*3+x*16+12],FIFO_7[256*3+x*16+12],FIFO_6[256*3+x*16+12],FIFO_5[256*3+x*16+12],FIFO_4[256*3+x*16+12],FIFO_3[256*3+x*16+12],FIFO_2[256*3+x*16+12],FIFO_1[256*3+x*16+12],FIFO_16[256*4+x*16+12],FIFO_15[256*4+x*16+12],FIFO_14[256*4+x*16+12],FIFO_13[256*4+x*16+12],FIFO_12[256*4+x*16+12],FIFO_11[256*4+x*16+12],FIFO_10[256*4+x*16+12],FIFO_9[256*4+x*16+12],FIFO_8[256*4+x*16+12],FIFO_7[256*4+x*16+12],FIFO_6[256*4+x*16+12],FIFO_5[256*4+x*16+12],FIFO_4[256*4+x*16+12],FIFO_3[256*4+x*16+12],FIFO_2[256*4+x*16+12],FIFO_1[256*4+x*16+12],FIFO_16[256*5+x*16+12],FIFO_15[256*5+x*16+12],FIFO_14[256*5+x*16+12],FIFO_13[256*5+x*16+12],FIFO_12[256*5+x*16+12],FIFO_11[256*5+x*16+12],FIFO_10[256*5+x*16+12],FIFO_9[256*5+x*16+12],FIFO_8[256*5+x*16+12],FIFO_7[256*5+x*16+12],FIFO_6[256*5+x*16+12],FIFO_5[256*5+x*16+12],FIFO_4[256*5+x*16+12],FIFO_3[256*5+x*16+12],FIFO_2[256*5+x*16+12],FIFO_1[256*5+x*16+12],FIFO_16[256*6+x*16+12],FIFO_15[256*6+x*16+12],FIFO_14[256*6+x*16+12],FIFO_13[256*6+x*16+12],FIFO_12[256*6+x*16+12],FIFO_11[256*6+x*16+12],FIFO_10[256*6+x*16+12],FIFO_9[256*6+x*16+12],FIFO_8[256*6+x*16+12],FIFO_7[256*6+x*16+12],FIFO_6[256*6+x*16+12],FIFO_5[256*6+x*16+12],FIFO_4[256*6+x*16+12],FIFO_3[256*6+x*16+12],FIFO_2[256*6+x*16+12],FIFO_1[256*6+x*16+12],FIFO_16[256*7+x*16+12],FIFO_15[256*7+x*16+12],FIFO_14[256*7+x*16+12],FIFO_13[256*7+x*16+12],FIFO_12[256*7+x*16+12],FIFO_11[256*7+x*16+12],FIFO_10[256*7+x*16+12],FIFO_9[256*7+x*16+12],FIFO_8[256*7+x*16+12],FIFO_7[256*7+x*16+12],FIFO_6[256*7+x*16+12],FIFO_5[256*7+x*16+12],FIFO_4[256*7+x*16+12],FIFO_3[256*7+x*16+12],FIFO_2[256*7+x*16+12],FIFO_1[256*7+x*16+12],FIFO_16[256*8+x*16+12],FIFO_15[256*8+x*16+12],FIFO_14[256*8+x*16+12],FIFO_13[256*8+x*16+12],FIFO_12[256*8+x*16+12],FIFO_11[256*8+x*16+12],FIFO_10[256*8+x*16+12],FIFO_9[256*8+x*16+12],FIFO_8[256*8+x*16+12],FIFO_7[256*8+x*16+12],FIFO_6[256*8+x*16+12],FIFO_5[256*8+x*16+12],FIFO_4[256*8+x*16+12],FIFO_3[256*8+x*16+12],FIFO_2[256*8+x*16+12],FIFO_1[256*8+x*16+12],FIFO_16[256*9+x*16+12],FIFO_15[256*9+x*16+12],FIFO_14[256*9+x*16+12],FIFO_13[256*9+x*16+12],FIFO_12[256*9+x*16+12],FIFO_11[256*9+x*16+12],FIFO_10[256*9+x*16+12],FIFO_9[256*9+x*16+12],FIFO_8[256*9+x*16+12],FIFO_7[256*9+x*16+12],FIFO_6[256*9+x*16+12],FIFO_5[256*9+x*16+12],FIFO_4[256*9+x*16+12],FIFO_3[256*9+x*16+12],FIFO_2[256*9+x*16+12],FIFO_1[256*9+x*16+12],FIFO_16[256*10+x*16+12],FIFO_15[256*10+x*16+12],FIFO_14[256*10+x*16+12],FIFO_13[256*10+x*16+12],FIFO_12[256*10+x*16+12],FIFO_11[256*10+x*16+12],FIFO_10[256*10+x*16+12],FIFO_9[256*10+x*16+12],FIFO_8[256*10+x*16+12],FIFO_7[256*10+x*16+12],FIFO_6[256*10+x*16+12],FIFO_5[256*10+x*16+12],FIFO_4[256*10+x*16+12],FIFO_3[256*10+x*16+12],FIFO_2[256*10+x*16+12],FIFO_1[256*10+x*16+12],FIFO_16[256*11+x*16+12],FIFO_15[256*11+x*16+12],FIFO_14[256*11+x*16+12],FIFO_13[256*11+x*16+12],FIFO_12[256*11+x*16+12],FIFO_11[256*11+x*16+12],FIFO_10[256*11+x*16+12],FIFO_9[256*11+x*16+12],FIFO_8[256*11+x*16+12],FIFO_7[256*11+x*16+12],FIFO_6[256*11+x*16+12],FIFO_5[256*11+x*16+12],FIFO_4[256*11+x*16+12],FIFO_3[256*11+x*16+12],FIFO_2[256*11+x*16+12],FIFO_1[256*11+x*16+12],FIFO_16[256*12+x*16+12],FIFO_15[256*12+x*16+12],FIFO_14[256*12+x*16+12],FIFO_13[256*12+x*16+12],FIFO_12[256*12+x*16+12],FIFO_11[256*12+x*16+12],FIFO_10[256*12+x*16+12],FIFO_9[256*12+x*16+12],FIFO_8[256*12+x*16+12],FIFO_7[256*12+x*16+12],FIFO_6[256*12+x*16+12],FIFO_5[256*12+x*16+12],FIFO_4[256*12+x*16+12],FIFO_3[256*12+x*16+12],FIFO_2[256*12+x*16+12],FIFO_1[256*12+x*16+12],FIFO_16[256*13+x*16+12],FIFO_15[256*13+x*16+12],FIFO_14[256*13+x*16+12],FIFO_13[256*13+x*16+12],FIFO_12[256*13+x*16+12],FIFO_11[256*13+x*16+12],FIFO_10[256*13+x*16+12],FIFO_9[256*13+x*16+12],FIFO_8[256*13+x*16+12],FIFO_7[256*13+x*16+12],FIFO_6[256*13+x*16+12],FIFO_5[256*13+x*16+12],FIFO_4[256*13+x*16+12],FIFO_3[256*13+x*16+12],FIFO_2[256*13+x*16+12],FIFO_1[256*13+x*16+12],FIFO_16[256*14+x*16+12],FIFO_15[256*14+x*16+12],FIFO_14[256*14+x*16+12],FIFO_13[256*14+x*16+12],FIFO_12[256*14+x*16+12],FIFO_11[256*14+x*16+12],FIFO_10[256*14+x*16+12],FIFO_9[256*14+x*16+12],FIFO_8[256*14+x*16+12],FIFO_7[256*14+x*16+12],FIFO_6[256*14+x*16+12],FIFO_5[256*14+x*16+12],FIFO_4[256*14+x*16+12],FIFO_3[256*14+x*16+12],FIFO_2[256*14+x*16+12],FIFO_1[256*14+x*16+12],FIFO_16[256*15+x*16+12],FIFO_15[256*15+x*16+12],FIFO_14[256*15+x*16+12],FIFO_13[256*15+x*16+12],FIFO_12[256*15+x*16+12],FIFO_11[256*15+x*16+12],FIFO_10[256*15+x*16+12],FIFO_9[256*15+x*16+12],FIFO_8[256*15+x*16+12],FIFO_7[256*15+x*16+12],FIFO_6[256*15+x*16+12],FIFO_5[256*15+x*16+12],FIFO_4[256*15+x*16+12],FIFO_3[256*15+x*16+12],FIFO_2[256*15+x*16+12],FIFO_1[256*15+x*16+12]}; 
                error_vector14 <= dec14 ^ {FIFO_16[256*0+x*16+13],FIFO_15[256*0+x*16+13],FIFO_14[256*0+x*16+13],FIFO_13[256*0+x*16+13],FIFO_12[256*0+x*16+13],FIFO_11[256*0+x*16+13],FIFO_10[256*0+x*16+13],FIFO_9[256*0+x*16+13],FIFO_8[256*0+x*16+13],FIFO_7[256*0+x*16+13],FIFO_6[256*0+x*16+13],FIFO_5[256*0+x*16+13],FIFO_4[256*0+x*16+13],FIFO_3[256*0+x*16+13],FIFO_2[256*0+x*16+13],FIFO_1[256*0+x*16+13],FIFO_16[256*1+x*16+13],FIFO_15[256*1+x*16+13],FIFO_14[256*1+x*16+13],FIFO_13[256*1+x*16+13],FIFO_12[256*1+x*16+13],FIFO_11[256*1+x*16+13],FIFO_10[256*1+x*16+13],FIFO_9[256*1+x*16+13],FIFO_8[256*1+x*16+13],FIFO_7[256*1+x*16+13],FIFO_6[256*1+x*16+13],FIFO_5[256*1+x*16+13],FIFO_4[256*1+x*16+13],FIFO_3[256*1+x*16+13],FIFO_2[256*1+x*16+13],FIFO_1[256*1+x*16+13],FIFO_16[256*2+x*16+13],FIFO_15[256*2+x*16+13],FIFO_14[256*2+x*16+13],FIFO_13[256*2+x*16+13],FIFO_12[256*2+x*16+13],FIFO_11[256*2+x*16+13],FIFO_10[256*2+x*16+13],FIFO_9[256*2+x*16+13],FIFO_8[256*2+x*16+13],FIFO_7[256*2+x*16+13],FIFO_6[256*2+x*16+13],FIFO_5[256*2+x*16+13],FIFO_4[256*2+x*16+13],FIFO_3[256*2+x*16+13],FIFO_2[256*2+x*16+13],FIFO_1[256*2+x*16+13],FIFO_16[256*3+x*16+13],FIFO_15[256*3+x*16+13],FIFO_14[256*3+x*16+13],FIFO_13[256*3+x*16+13],FIFO_12[256*3+x*16+13],FIFO_11[256*3+x*16+13],FIFO_10[256*3+x*16+13],FIFO_9[256*3+x*16+13],FIFO_8[256*3+x*16+13],FIFO_7[256*3+x*16+13],FIFO_6[256*3+x*16+13],FIFO_5[256*3+x*16+13],FIFO_4[256*3+x*16+13],FIFO_3[256*3+x*16+13],FIFO_2[256*3+x*16+13],FIFO_1[256*3+x*16+13],FIFO_16[256*4+x*16+13],FIFO_15[256*4+x*16+13],FIFO_14[256*4+x*16+13],FIFO_13[256*4+x*16+13],FIFO_12[256*4+x*16+13],FIFO_11[256*4+x*16+13],FIFO_10[256*4+x*16+13],FIFO_9[256*4+x*16+13],FIFO_8[256*4+x*16+13],FIFO_7[256*4+x*16+13],FIFO_6[256*4+x*16+13],FIFO_5[256*4+x*16+13],FIFO_4[256*4+x*16+13],FIFO_3[256*4+x*16+13],FIFO_2[256*4+x*16+13],FIFO_1[256*4+x*16+13],FIFO_16[256*5+x*16+13],FIFO_15[256*5+x*16+13],FIFO_14[256*5+x*16+13],FIFO_13[256*5+x*16+13],FIFO_12[256*5+x*16+13],FIFO_11[256*5+x*16+13],FIFO_10[256*5+x*16+13],FIFO_9[256*5+x*16+13],FIFO_8[256*5+x*16+13],FIFO_7[256*5+x*16+13],FIFO_6[256*5+x*16+13],FIFO_5[256*5+x*16+13],FIFO_4[256*5+x*16+13],FIFO_3[256*5+x*16+13],FIFO_2[256*5+x*16+13],FIFO_1[256*5+x*16+13],FIFO_16[256*6+x*16+13],FIFO_15[256*6+x*16+13],FIFO_14[256*6+x*16+13],FIFO_13[256*6+x*16+13],FIFO_12[256*6+x*16+13],FIFO_11[256*6+x*16+13],FIFO_10[256*6+x*16+13],FIFO_9[256*6+x*16+13],FIFO_8[256*6+x*16+13],FIFO_7[256*6+x*16+13],FIFO_6[256*6+x*16+13],FIFO_5[256*6+x*16+13],FIFO_4[256*6+x*16+13],FIFO_3[256*6+x*16+13],FIFO_2[256*6+x*16+13],FIFO_1[256*6+x*16+13],FIFO_16[256*7+x*16+13],FIFO_15[256*7+x*16+13],FIFO_14[256*7+x*16+13],FIFO_13[256*7+x*16+13],FIFO_12[256*7+x*16+13],FIFO_11[256*7+x*16+13],FIFO_10[256*7+x*16+13],FIFO_9[256*7+x*16+13],FIFO_8[256*7+x*16+13],FIFO_7[256*7+x*16+13],FIFO_6[256*7+x*16+13],FIFO_5[256*7+x*16+13],FIFO_4[256*7+x*16+13],FIFO_3[256*7+x*16+13],FIFO_2[256*7+x*16+13],FIFO_1[256*7+x*16+13],FIFO_16[256*8+x*16+13],FIFO_15[256*8+x*16+13],FIFO_14[256*8+x*16+13],FIFO_13[256*8+x*16+13],FIFO_12[256*8+x*16+13],FIFO_11[256*8+x*16+13],FIFO_10[256*8+x*16+13],FIFO_9[256*8+x*16+13],FIFO_8[256*8+x*16+13],FIFO_7[256*8+x*16+13],FIFO_6[256*8+x*16+13],FIFO_5[256*8+x*16+13],FIFO_4[256*8+x*16+13],FIFO_3[256*8+x*16+13],FIFO_2[256*8+x*16+13],FIFO_1[256*8+x*16+13],FIFO_16[256*9+x*16+13],FIFO_15[256*9+x*16+13],FIFO_14[256*9+x*16+13],FIFO_13[256*9+x*16+13],FIFO_12[256*9+x*16+13],FIFO_11[256*9+x*16+13],FIFO_10[256*9+x*16+13],FIFO_9[256*9+x*16+13],FIFO_8[256*9+x*16+13],FIFO_7[256*9+x*16+13],FIFO_6[256*9+x*16+13],FIFO_5[256*9+x*16+13],FIFO_4[256*9+x*16+13],FIFO_3[256*9+x*16+13],FIFO_2[256*9+x*16+13],FIFO_1[256*9+x*16+13],FIFO_16[256*10+x*16+13],FIFO_15[256*10+x*16+13],FIFO_14[256*10+x*16+13],FIFO_13[256*10+x*16+13],FIFO_12[256*10+x*16+13],FIFO_11[256*10+x*16+13],FIFO_10[256*10+x*16+13],FIFO_9[256*10+x*16+13],FIFO_8[256*10+x*16+13],FIFO_7[256*10+x*16+13],FIFO_6[256*10+x*16+13],FIFO_5[256*10+x*16+13],FIFO_4[256*10+x*16+13],FIFO_3[256*10+x*16+13],FIFO_2[256*10+x*16+13],FIFO_1[256*10+x*16+13],FIFO_16[256*11+x*16+13],FIFO_15[256*11+x*16+13],FIFO_14[256*11+x*16+13],FIFO_13[256*11+x*16+13],FIFO_12[256*11+x*16+13],FIFO_11[256*11+x*16+13],FIFO_10[256*11+x*16+13],FIFO_9[256*11+x*16+13],FIFO_8[256*11+x*16+13],FIFO_7[256*11+x*16+13],FIFO_6[256*11+x*16+13],FIFO_5[256*11+x*16+13],FIFO_4[256*11+x*16+13],FIFO_3[256*11+x*16+13],FIFO_2[256*11+x*16+13],FIFO_1[256*11+x*16+13],FIFO_16[256*12+x*16+13],FIFO_15[256*12+x*16+13],FIFO_14[256*12+x*16+13],FIFO_13[256*12+x*16+13],FIFO_12[256*12+x*16+13],FIFO_11[256*12+x*16+13],FIFO_10[256*12+x*16+13],FIFO_9[256*12+x*16+13],FIFO_8[256*12+x*16+13],FIFO_7[256*12+x*16+13],FIFO_6[256*12+x*16+13],FIFO_5[256*12+x*16+13],FIFO_4[256*12+x*16+13],FIFO_3[256*12+x*16+13],FIFO_2[256*12+x*16+13],FIFO_1[256*12+x*16+13],FIFO_16[256*13+x*16+13],FIFO_15[256*13+x*16+13],FIFO_14[256*13+x*16+13],FIFO_13[256*13+x*16+13],FIFO_12[256*13+x*16+13],FIFO_11[256*13+x*16+13],FIFO_10[256*13+x*16+13],FIFO_9[256*13+x*16+13],FIFO_8[256*13+x*16+13],FIFO_7[256*13+x*16+13],FIFO_6[256*13+x*16+13],FIFO_5[256*13+x*16+13],FIFO_4[256*13+x*16+13],FIFO_3[256*13+x*16+13],FIFO_2[256*13+x*16+13],FIFO_1[256*13+x*16+13],FIFO_16[256*14+x*16+13],FIFO_15[256*14+x*16+13],FIFO_14[256*14+x*16+13],FIFO_13[256*14+x*16+13],FIFO_12[256*14+x*16+13],FIFO_11[256*14+x*16+13],FIFO_10[256*14+x*16+13],FIFO_9[256*14+x*16+13],FIFO_8[256*14+x*16+13],FIFO_7[256*14+x*16+13],FIFO_6[256*14+x*16+13],FIFO_5[256*14+x*16+13],FIFO_4[256*14+x*16+13],FIFO_3[256*14+x*16+13],FIFO_2[256*14+x*16+13],FIFO_1[256*14+x*16+13],FIFO_16[256*15+x*16+13],FIFO_15[256*15+x*16+13],FIFO_14[256*15+x*16+13],FIFO_13[256*15+x*16+13],FIFO_12[256*15+x*16+13],FIFO_11[256*15+x*16+13],FIFO_10[256*15+x*16+13],FIFO_9[256*15+x*16+13],FIFO_8[256*15+x*16+13],FIFO_7[256*15+x*16+13],FIFO_6[256*15+x*16+13],FIFO_5[256*15+x*16+13],FIFO_4[256*15+x*16+13],FIFO_3[256*15+x*16+13],FIFO_2[256*15+x*16+13],FIFO_1[256*15+x*16+13]}; 
                error_vector15 <= dec15 ^ {FIFO_16[256*0+x*16+14],FIFO_15[256*0+x*16+14],FIFO_14[256*0+x*16+14],FIFO_13[256*0+x*16+14],FIFO_12[256*0+x*16+14],FIFO_11[256*0+x*16+14],FIFO_10[256*0+x*16+14],FIFO_9[256*0+x*16+14],FIFO_8[256*0+x*16+14],FIFO_7[256*0+x*16+14],FIFO_6[256*0+x*16+14],FIFO_5[256*0+x*16+14],FIFO_4[256*0+x*16+14],FIFO_3[256*0+x*16+14],FIFO_2[256*0+x*16+14],FIFO_1[256*0+x*16+14],FIFO_16[256*1+x*16+14],FIFO_15[256*1+x*16+14],FIFO_14[256*1+x*16+14],FIFO_13[256*1+x*16+14],FIFO_12[256*1+x*16+14],FIFO_11[256*1+x*16+14],FIFO_10[256*1+x*16+14],FIFO_9[256*1+x*16+14],FIFO_8[256*1+x*16+14],FIFO_7[256*1+x*16+14],FIFO_6[256*1+x*16+14],FIFO_5[256*1+x*16+14],FIFO_4[256*1+x*16+14],FIFO_3[256*1+x*16+14],FIFO_2[256*1+x*16+14],FIFO_1[256*1+x*16+14],FIFO_16[256*2+x*16+14],FIFO_15[256*2+x*16+14],FIFO_14[256*2+x*16+14],FIFO_13[256*2+x*16+14],FIFO_12[256*2+x*16+14],FIFO_11[256*2+x*16+14],FIFO_10[256*2+x*16+14],FIFO_9[256*2+x*16+14],FIFO_8[256*2+x*16+14],FIFO_7[256*2+x*16+14],FIFO_6[256*2+x*16+14],FIFO_5[256*2+x*16+14],FIFO_4[256*2+x*16+14],FIFO_3[256*2+x*16+14],FIFO_2[256*2+x*16+14],FIFO_1[256*2+x*16+14],FIFO_16[256*3+x*16+14],FIFO_15[256*3+x*16+14],FIFO_14[256*3+x*16+14],FIFO_13[256*3+x*16+14],FIFO_12[256*3+x*16+14],FIFO_11[256*3+x*16+14],FIFO_10[256*3+x*16+14],FIFO_9[256*3+x*16+14],FIFO_8[256*3+x*16+14],FIFO_7[256*3+x*16+14],FIFO_6[256*3+x*16+14],FIFO_5[256*3+x*16+14],FIFO_4[256*3+x*16+14],FIFO_3[256*3+x*16+14],FIFO_2[256*3+x*16+14],FIFO_1[256*3+x*16+14],FIFO_16[256*4+x*16+14],FIFO_15[256*4+x*16+14],FIFO_14[256*4+x*16+14],FIFO_13[256*4+x*16+14],FIFO_12[256*4+x*16+14],FIFO_11[256*4+x*16+14],FIFO_10[256*4+x*16+14],FIFO_9[256*4+x*16+14],FIFO_8[256*4+x*16+14],FIFO_7[256*4+x*16+14],FIFO_6[256*4+x*16+14],FIFO_5[256*4+x*16+14],FIFO_4[256*4+x*16+14],FIFO_3[256*4+x*16+14],FIFO_2[256*4+x*16+14],FIFO_1[256*4+x*16+14],FIFO_16[256*5+x*16+14],FIFO_15[256*5+x*16+14],FIFO_14[256*5+x*16+14],FIFO_13[256*5+x*16+14],FIFO_12[256*5+x*16+14],FIFO_11[256*5+x*16+14],FIFO_10[256*5+x*16+14],FIFO_9[256*5+x*16+14],FIFO_8[256*5+x*16+14],FIFO_7[256*5+x*16+14],FIFO_6[256*5+x*16+14],FIFO_5[256*5+x*16+14],FIFO_4[256*5+x*16+14],FIFO_3[256*5+x*16+14],FIFO_2[256*5+x*16+14],FIFO_1[256*5+x*16+14],FIFO_16[256*6+x*16+14],FIFO_15[256*6+x*16+14],FIFO_14[256*6+x*16+14],FIFO_13[256*6+x*16+14],FIFO_12[256*6+x*16+14],FIFO_11[256*6+x*16+14],FIFO_10[256*6+x*16+14],FIFO_9[256*6+x*16+14],FIFO_8[256*6+x*16+14],FIFO_7[256*6+x*16+14],FIFO_6[256*6+x*16+14],FIFO_5[256*6+x*16+14],FIFO_4[256*6+x*16+14],FIFO_3[256*6+x*16+14],FIFO_2[256*6+x*16+14],FIFO_1[256*6+x*16+14],FIFO_16[256*7+x*16+14],FIFO_15[256*7+x*16+14],FIFO_14[256*7+x*16+14],FIFO_13[256*7+x*16+14],FIFO_12[256*7+x*16+14],FIFO_11[256*7+x*16+14],FIFO_10[256*7+x*16+14],FIFO_9[256*7+x*16+14],FIFO_8[256*7+x*16+14],FIFO_7[256*7+x*16+14],FIFO_6[256*7+x*16+14],FIFO_5[256*7+x*16+14],FIFO_4[256*7+x*16+14],FIFO_3[256*7+x*16+14],FIFO_2[256*7+x*16+14],FIFO_1[256*7+x*16+14],FIFO_16[256*8+x*16+14],FIFO_15[256*8+x*16+14],FIFO_14[256*8+x*16+14],FIFO_13[256*8+x*16+14],FIFO_12[256*8+x*16+14],FIFO_11[256*8+x*16+14],FIFO_10[256*8+x*16+14],FIFO_9[256*8+x*16+14],FIFO_8[256*8+x*16+14],FIFO_7[256*8+x*16+14],FIFO_6[256*8+x*16+14],FIFO_5[256*8+x*16+14],FIFO_4[256*8+x*16+14],FIFO_3[256*8+x*16+14],FIFO_2[256*8+x*16+14],FIFO_1[256*8+x*16+14],FIFO_16[256*9+x*16+14],FIFO_15[256*9+x*16+14],FIFO_14[256*9+x*16+14],FIFO_13[256*9+x*16+14],FIFO_12[256*9+x*16+14],FIFO_11[256*9+x*16+14],FIFO_10[256*9+x*16+14],FIFO_9[256*9+x*16+14],FIFO_8[256*9+x*16+14],FIFO_7[256*9+x*16+14],FIFO_6[256*9+x*16+14],FIFO_5[256*9+x*16+14],FIFO_4[256*9+x*16+14],FIFO_3[256*9+x*16+14],FIFO_2[256*9+x*16+14],FIFO_1[256*9+x*16+14],FIFO_16[256*10+x*16+14],FIFO_15[256*10+x*16+14],FIFO_14[256*10+x*16+14],FIFO_13[256*10+x*16+14],FIFO_12[256*10+x*16+14],FIFO_11[256*10+x*16+14],FIFO_10[256*10+x*16+14],FIFO_9[256*10+x*16+14],FIFO_8[256*10+x*16+14],FIFO_7[256*10+x*16+14],FIFO_6[256*10+x*16+14],FIFO_5[256*10+x*16+14],FIFO_4[256*10+x*16+14],FIFO_3[256*10+x*16+14],FIFO_2[256*10+x*16+14],FIFO_1[256*10+x*16+14],FIFO_16[256*11+x*16+14],FIFO_15[256*11+x*16+14],FIFO_14[256*11+x*16+14],FIFO_13[256*11+x*16+14],FIFO_12[256*11+x*16+14],FIFO_11[256*11+x*16+14],FIFO_10[256*11+x*16+14],FIFO_9[256*11+x*16+14],FIFO_8[256*11+x*16+14],FIFO_7[256*11+x*16+14],FIFO_6[256*11+x*16+14],FIFO_5[256*11+x*16+14],FIFO_4[256*11+x*16+14],FIFO_3[256*11+x*16+14],FIFO_2[256*11+x*16+14],FIFO_1[256*11+x*16+14],FIFO_16[256*12+x*16+14],FIFO_15[256*12+x*16+14],FIFO_14[256*12+x*16+14],FIFO_13[256*12+x*16+14],FIFO_12[256*12+x*16+14],FIFO_11[256*12+x*16+14],FIFO_10[256*12+x*16+14],FIFO_9[256*12+x*16+14],FIFO_8[256*12+x*16+14],FIFO_7[256*12+x*16+14],FIFO_6[256*12+x*16+14],FIFO_5[256*12+x*16+14],FIFO_4[256*12+x*16+14],FIFO_3[256*12+x*16+14],FIFO_2[256*12+x*16+14],FIFO_1[256*12+x*16+14],FIFO_16[256*13+x*16+14],FIFO_15[256*13+x*16+14],FIFO_14[256*13+x*16+14],FIFO_13[256*13+x*16+14],FIFO_12[256*13+x*16+14],FIFO_11[256*13+x*16+14],FIFO_10[256*13+x*16+14],FIFO_9[256*13+x*16+14],FIFO_8[256*13+x*16+14],FIFO_7[256*13+x*16+14],FIFO_6[256*13+x*16+14],FIFO_5[256*13+x*16+14],FIFO_4[256*13+x*16+14],FIFO_3[256*13+x*16+14],FIFO_2[256*13+x*16+14],FIFO_1[256*13+x*16+14],FIFO_16[256*14+x*16+14],FIFO_15[256*14+x*16+14],FIFO_14[256*14+x*16+14],FIFO_13[256*14+x*16+14],FIFO_12[256*14+x*16+14],FIFO_11[256*14+x*16+14],FIFO_10[256*14+x*16+14],FIFO_9[256*14+x*16+14],FIFO_8[256*14+x*16+14],FIFO_7[256*14+x*16+14],FIFO_6[256*14+x*16+14],FIFO_5[256*14+x*16+14],FIFO_4[256*14+x*16+14],FIFO_3[256*14+x*16+14],FIFO_2[256*14+x*16+14],FIFO_1[256*14+x*16+14],FIFO_16[256*15+x*16+14],FIFO_15[256*15+x*16+14],FIFO_14[256*15+x*16+14],FIFO_13[256*15+x*16+14],FIFO_12[256*15+x*16+14],FIFO_11[256*15+x*16+14],FIFO_10[256*15+x*16+14],FIFO_9[256*15+x*16+14],FIFO_8[256*15+x*16+14],FIFO_7[256*15+x*16+14],FIFO_6[256*15+x*16+14],FIFO_5[256*15+x*16+14],FIFO_4[256*15+x*16+14],FIFO_3[256*15+x*16+14],FIFO_2[256*15+x*16+14],FIFO_1[256*15+x*16+14]}; 
                error_vector16 <= dec16 ^ {FIFO_16[256*0+x*16+15],FIFO_15[256*0+x*16+15],FIFO_14[256*0+x*16+15],FIFO_13[256*0+x*16+15],FIFO_12[256*0+x*16+15],FIFO_11[256*0+x*16+15],FIFO_10[256*0+x*16+15],FIFO_9[256*0+x*16+15],FIFO_8[256*0+x*16+15],FIFO_7[256*0+x*16+15],FIFO_6[256*0+x*16+15],FIFO_5[256*0+x*16+15],FIFO_4[256*0+x*16+15],FIFO_3[256*0+x*16+15],FIFO_2[256*0+x*16+15],FIFO_1[256*0+x*16+15],FIFO_16[256*1+x*16+15],FIFO_15[256*1+x*16+15],FIFO_14[256*1+x*16+15],FIFO_13[256*1+x*16+15],FIFO_12[256*1+x*16+15],FIFO_11[256*1+x*16+15],FIFO_10[256*1+x*16+15],FIFO_9[256*1+x*16+15],FIFO_8[256*1+x*16+15],FIFO_7[256*1+x*16+15],FIFO_6[256*1+x*16+15],FIFO_5[256*1+x*16+15],FIFO_4[256*1+x*16+15],FIFO_3[256*1+x*16+15],FIFO_2[256*1+x*16+15],FIFO_1[256*1+x*16+15],FIFO_16[256*2+x*16+15],FIFO_15[256*2+x*16+15],FIFO_14[256*2+x*16+15],FIFO_13[256*2+x*16+15],FIFO_12[256*2+x*16+15],FIFO_11[256*2+x*16+15],FIFO_10[256*2+x*16+15],FIFO_9[256*2+x*16+15],FIFO_8[256*2+x*16+15],FIFO_7[256*2+x*16+15],FIFO_6[256*2+x*16+15],FIFO_5[256*2+x*16+15],FIFO_4[256*2+x*16+15],FIFO_3[256*2+x*16+15],FIFO_2[256*2+x*16+15],FIFO_1[256*2+x*16+15],FIFO_16[256*3+x*16+15],FIFO_15[256*3+x*16+15],FIFO_14[256*3+x*16+15],FIFO_13[256*3+x*16+15],FIFO_12[256*3+x*16+15],FIFO_11[256*3+x*16+15],FIFO_10[256*3+x*16+15],FIFO_9[256*3+x*16+15],FIFO_8[256*3+x*16+15],FIFO_7[256*3+x*16+15],FIFO_6[256*3+x*16+15],FIFO_5[256*3+x*16+15],FIFO_4[256*3+x*16+15],FIFO_3[256*3+x*16+15],FIFO_2[256*3+x*16+15],FIFO_1[256*3+x*16+15],FIFO_16[256*4+x*16+15],FIFO_15[256*4+x*16+15],FIFO_14[256*4+x*16+15],FIFO_13[256*4+x*16+15],FIFO_12[256*4+x*16+15],FIFO_11[256*4+x*16+15],FIFO_10[256*4+x*16+15],FIFO_9[256*4+x*16+15],FIFO_8[256*4+x*16+15],FIFO_7[256*4+x*16+15],FIFO_6[256*4+x*16+15],FIFO_5[256*4+x*16+15],FIFO_4[256*4+x*16+15],FIFO_3[256*4+x*16+15],FIFO_2[256*4+x*16+15],FIFO_1[256*4+x*16+15],FIFO_16[256*5+x*16+15],FIFO_15[256*5+x*16+15],FIFO_14[256*5+x*16+15],FIFO_13[256*5+x*16+15],FIFO_12[256*5+x*16+15],FIFO_11[256*5+x*16+15],FIFO_10[256*5+x*16+15],FIFO_9[256*5+x*16+15],FIFO_8[256*5+x*16+15],FIFO_7[256*5+x*16+15],FIFO_6[256*5+x*16+15],FIFO_5[256*5+x*16+15],FIFO_4[256*5+x*16+15],FIFO_3[256*5+x*16+15],FIFO_2[256*5+x*16+15],FIFO_1[256*5+x*16+15],FIFO_16[256*6+x*16+15],FIFO_15[256*6+x*16+15],FIFO_14[256*6+x*16+15],FIFO_13[256*6+x*16+15],FIFO_12[256*6+x*16+15],FIFO_11[256*6+x*16+15],FIFO_10[256*6+x*16+15],FIFO_9[256*6+x*16+15],FIFO_8[256*6+x*16+15],FIFO_7[256*6+x*16+15],FIFO_6[256*6+x*16+15],FIFO_5[256*6+x*16+15],FIFO_4[256*6+x*16+15],FIFO_3[256*6+x*16+15],FIFO_2[256*6+x*16+15],FIFO_1[256*6+x*16+15],FIFO_16[256*7+x*16+15],FIFO_15[256*7+x*16+15],FIFO_14[256*7+x*16+15],FIFO_13[256*7+x*16+15],FIFO_12[256*7+x*16+15],FIFO_11[256*7+x*16+15],FIFO_10[256*7+x*16+15],FIFO_9[256*7+x*16+15],FIFO_8[256*7+x*16+15],FIFO_7[256*7+x*16+15],FIFO_6[256*7+x*16+15],FIFO_5[256*7+x*16+15],FIFO_4[256*7+x*16+15],FIFO_3[256*7+x*16+15],FIFO_2[256*7+x*16+15],FIFO_1[256*7+x*16+15],FIFO_16[256*8+x*16+15],FIFO_15[256*8+x*16+15],FIFO_14[256*8+x*16+15],FIFO_13[256*8+x*16+15],FIFO_12[256*8+x*16+15],FIFO_11[256*8+x*16+15],FIFO_10[256*8+x*16+15],FIFO_9[256*8+x*16+15],FIFO_8[256*8+x*16+15],FIFO_7[256*8+x*16+15],FIFO_6[256*8+x*16+15],FIFO_5[256*8+x*16+15],FIFO_4[256*8+x*16+15],FIFO_3[256*8+x*16+15],FIFO_2[256*8+x*16+15],FIFO_1[256*8+x*16+15],FIFO_16[256*9+x*16+15],FIFO_15[256*9+x*16+15],FIFO_14[256*9+x*16+15],FIFO_13[256*9+x*16+15],FIFO_12[256*9+x*16+15],FIFO_11[256*9+x*16+15],FIFO_10[256*9+x*16+15],FIFO_9[256*9+x*16+15],FIFO_8[256*9+x*16+15],FIFO_7[256*9+x*16+15],FIFO_6[256*9+x*16+15],FIFO_5[256*9+x*16+15],FIFO_4[256*9+x*16+15],FIFO_3[256*9+x*16+15],FIFO_2[256*9+x*16+15],FIFO_1[256*9+x*16+15],FIFO_16[256*10+x*16+15],FIFO_15[256*10+x*16+15],FIFO_14[256*10+x*16+15],FIFO_13[256*10+x*16+15],FIFO_12[256*10+x*16+15],FIFO_11[256*10+x*16+15],FIFO_10[256*10+x*16+15],FIFO_9[256*10+x*16+15],FIFO_8[256*10+x*16+15],FIFO_7[256*10+x*16+15],FIFO_6[256*10+x*16+15],FIFO_5[256*10+x*16+15],FIFO_4[256*10+x*16+15],FIFO_3[256*10+x*16+15],FIFO_2[256*10+x*16+15],FIFO_1[256*10+x*16+15],FIFO_16[256*11+x*16+15],FIFO_15[256*11+x*16+15],FIFO_14[256*11+x*16+15],FIFO_13[256*11+x*16+15],FIFO_12[256*11+x*16+15],FIFO_11[256*11+x*16+15],FIFO_10[256*11+x*16+15],FIFO_9[256*11+x*16+15],FIFO_8[256*11+x*16+15],FIFO_7[256*11+x*16+15],FIFO_6[256*11+x*16+15],FIFO_5[256*11+x*16+15],FIFO_4[256*11+x*16+15],FIFO_3[256*11+x*16+15],FIFO_2[256*11+x*16+15],FIFO_1[256*11+x*16+15],FIFO_16[256*12+x*16+15],FIFO_15[256*12+x*16+15],FIFO_14[256*12+x*16+15],FIFO_13[256*12+x*16+15],FIFO_12[256*12+x*16+15],FIFO_11[256*12+x*16+15],FIFO_10[256*12+x*16+15],FIFO_9[256*12+x*16+15],FIFO_8[256*12+x*16+15],FIFO_7[256*12+x*16+15],FIFO_6[256*12+x*16+15],FIFO_5[256*12+x*16+15],FIFO_4[256*12+x*16+15],FIFO_3[256*12+x*16+15],FIFO_2[256*12+x*16+15],FIFO_1[256*12+x*16+15],FIFO_16[256*13+x*16+15],FIFO_15[256*13+x*16+15],FIFO_14[256*13+x*16+15],FIFO_13[256*13+x*16+15],FIFO_12[256*13+x*16+15],FIFO_11[256*13+x*16+15],FIFO_10[256*13+x*16+15],FIFO_9[256*13+x*16+15],FIFO_8[256*13+x*16+15],FIFO_7[256*13+x*16+15],FIFO_6[256*13+x*16+15],FIFO_5[256*13+x*16+15],FIFO_4[256*13+x*16+15],FIFO_3[256*13+x*16+15],FIFO_2[256*13+x*16+15],FIFO_1[256*13+x*16+15],FIFO_16[256*14+x*16+15],FIFO_15[256*14+x*16+15],FIFO_14[256*14+x*16+15],FIFO_13[256*14+x*16+15],FIFO_12[256*14+x*16+15],FIFO_11[256*14+x*16+15],FIFO_10[256*14+x*16+15],FIFO_9[256*14+x*16+15],FIFO_8[256*14+x*16+15],FIFO_7[256*14+x*16+15],FIFO_6[256*14+x*16+15],FIFO_5[256*14+x*16+15],FIFO_4[256*14+x*16+15],FIFO_3[256*14+x*16+15],FIFO_2[256*14+x*16+15],FIFO_1[256*14+x*16+15],FIFO_16[256*15+x*16+15],FIFO_15[256*15+x*16+15],FIFO_14[256*15+x*16+15],FIFO_13[256*15+x*16+15],FIFO_12[256*15+x*16+15],FIFO_11[256*15+x*16+15],FIFO_10[256*15+x*16+15],FIFO_9[256*15+x*16+15],FIFO_8[256*15+x*16+15],FIFO_7[256*15+x*16+15],FIFO_6[256*15+x*16+15],FIFO_5[256*15+x*16+15],FIFO_4[256*15+x*16+15],FIFO_3[256*15+x*16+15],FIFO_2[256*15+x*16+15],FIFO_1[256*15+x*16+15]}; 
            
            end else begin
                x <= 5'b0;
                
                error_vector1 <= 0;
                error_vector2 <= 0;
                error_vector3 <= 0;
                error_vector4 <= 0;
                error_vector5 <= 0;
                error_vector6 <= 0;
                error_vector7 <= 0;
                error_vector8 <= 0;
                error_vector9 <= 0;
                error_vector10 <= 0;
                error_vector11 <= 0;
                error_vector12 <= 0;
                error_vector13 <= 0;
                error_vector14 <= 0;
                error_vector15 <= 0;
                error_vector16 <= 0;
            end

            errs1_u <= error_u_vector1[0] + error_u_vector1[1] + error_u_vector1[2] + error_u_vector1[3] + error_u_vector1[4] + error_u_vector1[5] + error_u_vector1[6] + error_u_vector1[7] + error_u_vector1[8] + error_u_vector1[9] + error_u_vector1[10] + error_u_vector1[11] + error_u_vector1[12] + error_u_vector1[13] + error_u_vector1[14] + error_u_vector1[15] + error_u_vector1[16] + error_u_vector1[17] + error_u_vector1[18] + error_u_vector1[19] + error_u_vector1[20] + error_u_vector1[21] + error_u_vector1[22] + error_u_vector1[23] + error_u_vector1[24] + error_u_vector1[25] + error_u_vector1[26] + error_u_vector1[27] + error_u_vector1[28] + error_u_vector1[29] + error_u_vector1[30] + error_u_vector1[31] + error_u_vector1[32] + error_u_vector1[33] + error_u_vector1[34] + error_u_vector1[35] + error_u_vector1[36] + error_u_vector1[37] + error_u_vector1[38] + error_u_vector1[39] + error_u_vector1[40] + error_u_vector1[41] + error_u_vector1[42] + error_u_vector1[43] + error_u_vector1[44] + error_u_vector1[45] + error_u_vector1[46] + error_u_vector1[47] + error_u_vector1[48] + error_u_vector1[49] + error_u_vector1[50] + error_u_vector1[51] + error_u_vector1[52] + error_u_vector1[53] + error_u_vector1[54] + error_u_vector1[55] + error_u_vector1[56] + error_u_vector1[57] + error_u_vector1[58] + error_u_vector1[59] + error_u_vector1[60] + error_u_vector1[61] + error_u_vector1[62] + error_u_vector1[63] + error_u_vector1[64] + error_u_vector1[65] + error_u_vector1[66] + error_u_vector1[67] + error_u_vector1[68] + error_u_vector1[69] + error_u_vector1[70] + error_u_vector1[71] + error_u_vector1[72] + error_u_vector1[73] + error_u_vector1[74] + error_u_vector1[75] + error_u_vector1[76] + error_u_vector1[77] + error_u_vector1[78] + error_u_vector1[79] + error_u_vector1[80] + error_u_vector1[81] + error_u_vector1[82] + error_u_vector1[83] + error_u_vector1[84] + error_u_vector1[85] + error_u_vector1[86] + error_u_vector1[87] + error_u_vector1[88] + error_u_vector1[89] + error_u_vector1[90] + error_u_vector1[91] + error_u_vector1[92] + error_u_vector1[93] + error_u_vector1[94] + error_u_vector1[95] + error_u_vector1[96] + error_u_vector1[97] + error_u_vector1[98] + error_u_vector1[99] + error_u_vector1[100] + error_u_vector1[101] + error_u_vector1[102] + error_u_vector1[103] + error_u_vector1[104] + error_u_vector1[105] + error_u_vector1[106] + error_u_vector1[107] + error_u_vector1[108] + error_u_vector1[109] + error_u_vector1[110] + error_u_vector1[111] + error_u_vector1[112] + error_u_vector1[113] + error_u_vector1[114] + error_u_vector1[115] + error_u_vector1[116] + error_u_vector1[117] + error_u_vector1[118] + error_u_vector1[119] + error_u_vector1[120] + error_u_vector1[121] + error_u_vector1[122] + error_u_vector1[123] + error_u_vector1[124] + error_u_vector1[125] + error_u_vector1[126] + error_u_vector1[127] + error_u_vector1[128] + error_u_vector1[129] + error_u_vector1[130] + error_u_vector1[131] + error_u_vector1[132] + error_u_vector1[133] + error_u_vector1[134] + error_u_vector1[135] + error_u_vector1[136] + error_u_vector1[137] + error_u_vector1[138] + error_u_vector1[139] + error_u_vector1[140] + error_u_vector1[141] + error_u_vector1[142] + error_u_vector1[143] + error_u_vector1[144] + error_u_vector1[145] + error_u_vector1[146] + error_u_vector1[147] + error_u_vector1[148] + error_u_vector1[149] + error_u_vector1[150] + error_u_vector1[151] + error_u_vector1[152] + error_u_vector1[153] + error_u_vector1[154] + error_u_vector1[155] + error_u_vector1[156] + error_u_vector1[157] + error_u_vector1[158] + error_u_vector1[159] + error_u_vector1[160] + error_u_vector1[161] + error_u_vector1[162] + error_u_vector1[163] + error_u_vector1[164] + error_u_vector1[165] + error_u_vector1[166] + error_u_vector1[167] + error_u_vector1[168] + error_u_vector1[169] + error_u_vector1[170] + error_u_vector1[171] + error_u_vector1[172] + error_u_vector1[173] + error_u_vector1[174] + error_u_vector1[175] + error_u_vector1[176] + error_u_vector1[177] + error_u_vector1[178] + error_u_vector1[179] + error_u_vector1[180] + error_u_vector1[181] + error_u_vector1[182] + error_u_vector1[183] + error_u_vector1[184] + error_u_vector1[185] + error_u_vector1[186] + error_u_vector1[187] + error_u_vector1[188] + error_u_vector1[189] + error_u_vector1[190] + error_u_vector1[191] + error_u_vector1[192] + error_u_vector1[193] + error_u_vector1[194] + error_u_vector1[195] + error_u_vector1[196] + error_u_vector1[197] + error_u_vector1[198] + error_u_vector1[199] + error_u_vector1[200] + error_u_vector1[201] + error_u_vector1[202] + error_u_vector1[203] + error_u_vector1[204] + error_u_vector1[205] + error_u_vector1[206] + error_u_vector1[207] + error_u_vector1[208] + error_u_vector1[209] + error_u_vector1[210] + error_u_vector1[211] + error_u_vector1[212] + error_u_vector1[213] + error_u_vector1[214] + error_u_vector1[215] + error_u_vector1[216] + error_u_vector1[217] + error_u_vector1[218] + error_u_vector1[219] + error_u_vector1[220] + error_u_vector1[221] + error_u_vector1[222] + error_u_vector1[223] + error_u_vector1[224] + error_u_vector1[225] + error_u_vector1[226] + error_u_vector1[227] + error_u_vector1[228] + error_u_vector1[229] + error_u_vector1[230] + error_u_vector1[231] + error_u_vector1[232] + error_u_vector1[233] + error_u_vector1[234] + error_u_vector1[235] + error_u_vector1[236] + error_u_vector1[237] + error_u_vector1[238]; 
            errs2_u <= error_u_vector2[0] + error_u_vector2[1] + error_u_vector2[2] + error_u_vector2[3] + error_u_vector2[4] + error_u_vector2[5] + error_u_vector2[6] + error_u_vector2[7] + error_u_vector2[8] + error_u_vector2[9] + error_u_vector2[10] + error_u_vector2[11] + error_u_vector2[12] + error_u_vector2[13] + error_u_vector2[14] + error_u_vector2[15] + error_u_vector2[16] + error_u_vector2[17] + error_u_vector2[18] + error_u_vector2[19] + error_u_vector2[20] + error_u_vector2[21] + error_u_vector2[22] + error_u_vector2[23] + error_u_vector2[24] + error_u_vector2[25] + error_u_vector2[26] + error_u_vector2[27] + error_u_vector2[28] + error_u_vector2[29] + error_u_vector2[30] + error_u_vector2[31] + error_u_vector2[32] + error_u_vector2[33] + error_u_vector2[34] + error_u_vector2[35] + error_u_vector2[36] + error_u_vector2[37] + error_u_vector2[38] + error_u_vector2[39] + error_u_vector2[40] + error_u_vector2[41] + error_u_vector2[42] + error_u_vector2[43] + error_u_vector2[44] + error_u_vector2[45] + error_u_vector2[46] + error_u_vector2[47] + error_u_vector2[48] + error_u_vector2[49] + error_u_vector2[50] + error_u_vector2[51] + error_u_vector2[52] + error_u_vector2[53] + error_u_vector2[54] + error_u_vector2[55] + error_u_vector2[56] + error_u_vector2[57] + error_u_vector2[58] + error_u_vector2[59] + error_u_vector2[60] + error_u_vector2[61] + error_u_vector2[62] + error_u_vector2[63] + error_u_vector2[64] + error_u_vector2[65] + error_u_vector2[66] + error_u_vector2[67] + error_u_vector2[68] + error_u_vector2[69] + error_u_vector2[70] + error_u_vector2[71] + error_u_vector2[72] + error_u_vector2[73] + error_u_vector2[74] + error_u_vector2[75] + error_u_vector2[76] + error_u_vector2[77] + error_u_vector2[78] + error_u_vector2[79] + error_u_vector2[80] + error_u_vector2[81] + error_u_vector2[82] + error_u_vector2[83] + error_u_vector2[84] + error_u_vector2[85] + error_u_vector2[86] + error_u_vector2[87] + error_u_vector2[88] + error_u_vector2[89] + error_u_vector2[90] + error_u_vector2[91] + error_u_vector2[92] + error_u_vector2[93] + error_u_vector2[94] + error_u_vector2[95] + error_u_vector2[96] + error_u_vector2[97] + error_u_vector2[98] + error_u_vector2[99] + error_u_vector2[100] + error_u_vector2[101] + error_u_vector2[102] + error_u_vector2[103] + error_u_vector2[104] + error_u_vector2[105] + error_u_vector2[106] + error_u_vector2[107] + error_u_vector2[108] + error_u_vector2[109] + error_u_vector2[110] + error_u_vector2[111] + error_u_vector2[112] + error_u_vector2[113] + error_u_vector2[114] + error_u_vector2[115] + error_u_vector2[116] + error_u_vector2[117] + error_u_vector2[118] + error_u_vector2[119] + error_u_vector2[120] + error_u_vector2[121] + error_u_vector2[122] + error_u_vector2[123] + error_u_vector2[124] + error_u_vector2[125] + error_u_vector2[126] + error_u_vector2[127] + error_u_vector2[128] + error_u_vector2[129] + error_u_vector2[130] + error_u_vector2[131] + error_u_vector2[132] + error_u_vector2[133] + error_u_vector2[134] + error_u_vector2[135] + error_u_vector2[136] + error_u_vector2[137] + error_u_vector2[138] + error_u_vector2[139] + error_u_vector2[140] + error_u_vector2[141] + error_u_vector2[142] + error_u_vector2[143] + error_u_vector2[144] + error_u_vector2[145] + error_u_vector2[146] + error_u_vector2[147] + error_u_vector2[148] + error_u_vector2[149] + error_u_vector2[150] + error_u_vector2[151] + error_u_vector2[152] + error_u_vector2[153] + error_u_vector2[154] + error_u_vector2[155] + error_u_vector2[156] + error_u_vector2[157] + error_u_vector2[158] + error_u_vector2[159] + error_u_vector2[160] + error_u_vector2[161] + error_u_vector2[162] + error_u_vector2[163] + error_u_vector2[164] + error_u_vector2[165] + error_u_vector2[166] + error_u_vector2[167] + error_u_vector2[168] + error_u_vector2[169] + error_u_vector2[170] + error_u_vector2[171] + error_u_vector2[172] + error_u_vector2[173] + error_u_vector2[174] + error_u_vector2[175] + error_u_vector2[176] + error_u_vector2[177] + error_u_vector2[178] + error_u_vector2[179] + error_u_vector2[180] + error_u_vector2[181] + error_u_vector2[182] + error_u_vector2[183] + error_u_vector2[184] + error_u_vector2[185] + error_u_vector2[186] + error_u_vector2[187] + error_u_vector2[188] + error_u_vector2[189] + error_u_vector2[190] + error_u_vector2[191] + error_u_vector2[192] + error_u_vector2[193] + error_u_vector2[194] + error_u_vector2[195] + error_u_vector2[196] + error_u_vector2[197] + error_u_vector2[198] + error_u_vector2[199] + error_u_vector2[200] + error_u_vector2[201] + error_u_vector2[202] + error_u_vector2[203] + error_u_vector2[204] + error_u_vector2[205] + error_u_vector2[206] + error_u_vector2[207] + error_u_vector2[208] + error_u_vector2[209] + error_u_vector2[210] + error_u_vector2[211] + error_u_vector2[212] + error_u_vector2[213] + error_u_vector2[214] + error_u_vector2[215] + error_u_vector2[216] + error_u_vector2[217] + error_u_vector2[218] + error_u_vector2[219] + error_u_vector2[220] + error_u_vector2[221] + error_u_vector2[222] + error_u_vector2[223] + error_u_vector2[224] + error_u_vector2[225] + error_u_vector2[226] + error_u_vector2[227] + error_u_vector2[228] + error_u_vector2[229] + error_u_vector2[230] + error_u_vector2[231] + error_u_vector2[232] + error_u_vector2[233] + error_u_vector2[234] + error_u_vector2[235] + error_u_vector2[236] + error_u_vector2[237] + error_u_vector2[238]; 
            errs3_u <= error_u_vector3[0] + error_u_vector3[1] + error_u_vector3[2] + error_u_vector3[3] + error_u_vector3[4] + error_u_vector3[5] + error_u_vector3[6] + error_u_vector3[7] + error_u_vector3[8] + error_u_vector3[9] + error_u_vector3[10] + error_u_vector3[11] + error_u_vector3[12] + error_u_vector3[13] + error_u_vector3[14] + error_u_vector3[15] + error_u_vector3[16] + error_u_vector3[17] + error_u_vector3[18] + error_u_vector3[19] + error_u_vector3[20] + error_u_vector3[21] + error_u_vector3[22] + error_u_vector3[23] + error_u_vector3[24] + error_u_vector3[25] + error_u_vector3[26] + error_u_vector3[27] + error_u_vector3[28] + error_u_vector3[29] + error_u_vector3[30] + error_u_vector3[31] + error_u_vector3[32] + error_u_vector3[33] + error_u_vector3[34] + error_u_vector3[35] + error_u_vector3[36] + error_u_vector3[37] + error_u_vector3[38] + error_u_vector3[39] + error_u_vector3[40] + error_u_vector3[41] + error_u_vector3[42] + error_u_vector3[43] + error_u_vector3[44] + error_u_vector3[45] + error_u_vector3[46] + error_u_vector3[47] + error_u_vector3[48] + error_u_vector3[49] + error_u_vector3[50] + error_u_vector3[51] + error_u_vector3[52] + error_u_vector3[53] + error_u_vector3[54] + error_u_vector3[55] + error_u_vector3[56] + error_u_vector3[57] + error_u_vector3[58] + error_u_vector3[59] + error_u_vector3[60] + error_u_vector3[61] + error_u_vector3[62] + error_u_vector3[63] + error_u_vector3[64] + error_u_vector3[65] + error_u_vector3[66] + error_u_vector3[67] + error_u_vector3[68] + error_u_vector3[69] + error_u_vector3[70] + error_u_vector3[71] + error_u_vector3[72] + error_u_vector3[73] + error_u_vector3[74] + error_u_vector3[75] + error_u_vector3[76] + error_u_vector3[77] + error_u_vector3[78] + error_u_vector3[79] + error_u_vector3[80] + error_u_vector3[81] + error_u_vector3[82] + error_u_vector3[83] + error_u_vector3[84] + error_u_vector3[85] + error_u_vector3[86] + error_u_vector3[87] + error_u_vector3[88] + error_u_vector3[89] + error_u_vector3[90] + error_u_vector3[91] + error_u_vector3[92] + error_u_vector3[93] + error_u_vector3[94] + error_u_vector3[95] + error_u_vector3[96] + error_u_vector3[97] + error_u_vector3[98] + error_u_vector3[99] + error_u_vector3[100] + error_u_vector3[101] + error_u_vector3[102] + error_u_vector3[103] + error_u_vector3[104] + error_u_vector3[105] + error_u_vector3[106] + error_u_vector3[107] + error_u_vector3[108] + error_u_vector3[109] + error_u_vector3[110] + error_u_vector3[111] + error_u_vector3[112] + error_u_vector3[113] + error_u_vector3[114] + error_u_vector3[115] + error_u_vector3[116] + error_u_vector3[117] + error_u_vector3[118] + error_u_vector3[119] + error_u_vector3[120] + error_u_vector3[121] + error_u_vector3[122] + error_u_vector3[123] + error_u_vector3[124] + error_u_vector3[125] + error_u_vector3[126] + error_u_vector3[127] + error_u_vector3[128] + error_u_vector3[129] + error_u_vector3[130] + error_u_vector3[131] + error_u_vector3[132] + error_u_vector3[133] + error_u_vector3[134] + error_u_vector3[135] + error_u_vector3[136] + error_u_vector3[137] + error_u_vector3[138] + error_u_vector3[139] + error_u_vector3[140] + error_u_vector3[141] + error_u_vector3[142] + error_u_vector3[143] + error_u_vector3[144] + error_u_vector3[145] + error_u_vector3[146] + error_u_vector3[147] + error_u_vector3[148] + error_u_vector3[149] + error_u_vector3[150] + error_u_vector3[151] + error_u_vector3[152] + error_u_vector3[153] + error_u_vector3[154] + error_u_vector3[155] + error_u_vector3[156] + error_u_vector3[157] + error_u_vector3[158] + error_u_vector3[159] + error_u_vector3[160] + error_u_vector3[161] + error_u_vector3[162] + error_u_vector3[163] + error_u_vector3[164] + error_u_vector3[165] + error_u_vector3[166] + error_u_vector3[167] + error_u_vector3[168] + error_u_vector3[169] + error_u_vector3[170] + error_u_vector3[171] + error_u_vector3[172] + error_u_vector3[173] + error_u_vector3[174] + error_u_vector3[175] + error_u_vector3[176] + error_u_vector3[177] + error_u_vector3[178] + error_u_vector3[179] + error_u_vector3[180] + error_u_vector3[181] + error_u_vector3[182] + error_u_vector3[183] + error_u_vector3[184] + error_u_vector3[185] + error_u_vector3[186] + error_u_vector3[187] + error_u_vector3[188] + error_u_vector3[189] + error_u_vector3[190] + error_u_vector3[191] + error_u_vector3[192] + error_u_vector3[193] + error_u_vector3[194] + error_u_vector3[195] + error_u_vector3[196] + error_u_vector3[197] + error_u_vector3[198] + error_u_vector3[199] + error_u_vector3[200] + error_u_vector3[201] + error_u_vector3[202] + error_u_vector3[203] + error_u_vector3[204] + error_u_vector3[205] + error_u_vector3[206] + error_u_vector3[207] + error_u_vector3[208] + error_u_vector3[209] + error_u_vector3[210] + error_u_vector3[211] + error_u_vector3[212] + error_u_vector3[213] + error_u_vector3[214] + error_u_vector3[215] + error_u_vector3[216] + error_u_vector3[217] + error_u_vector3[218] + error_u_vector3[219] + error_u_vector3[220] + error_u_vector3[221] + error_u_vector3[222] + error_u_vector3[223] + error_u_vector3[224] + error_u_vector3[225] + error_u_vector3[226] + error_u_vector3[227] + error_u_vector3[228] + error_u_vector3[229] + error_u_vector3[230] + error_u_vector3[231] + error_u_vector3[232] + error_u_vector3[233] + error_u_vector3[234] + error_u_vector3[235] + error_u_vector3[236] + error_u_vector3[237] + error_u_vector3[238]; 
            errs4_u <= error_u_vector4[0] + error_u_vector4[1] + error_u_vector4[2] + error_u_vector4[3] + error_u_vector4[4] + error_u_vector4[5] + error_u_vector4[6] + error_u_vector4[7] + error_u_vector4[8] + error_u_vector4[9] + error_u_vector4[10] + error_u_vector4[11] + error_u_vector4[12] + error_u_vector4[13] + error_u_vector4[14] + error_u_vector4[15] + error_u_vector4[16] + error_u_vector4[17] + error_u_vector4[18] + error_u_vector4[19] + error_u_vector4[20] + error_u_vector4[21] + error_u_vector4[22] + error_u_vector4[23] + error_u_vector4[24] + error_u_vector4[25] + error_u_vector4[26] + error_u_vector4[27] + error_u_vector4[28] + error_u_vector4[29] + error_u_vector4[30] + error_u_vector4[31] + error_u_vector4[32] + error_u_vector4[33] + error_u_vector4[34] + error_u_vector4[35] + error_u_vector4[36] + error_u_vector4[37] + error_u_vector4[38] + error_u_vector4[39] + error_u_vector4[40] + error_u_vector4[41] + error_u_vector4[42] + error_u_vector4[43] + error_u_vector4[44] + error_u_vector4[45] + error_u_vector4[46] + error_u_vector4[47] + error_u_vector4[48] + error_u_vector4[49] + error_u_vector4[50] + error_u_vector4[51] + error_u_vector4[52] + error_u_vector4[53] + error_u_vector4[54] + error_u_vector4[55] + error_u_vector4[56] + error_u_vector4[57] + error_u_vector4[58] + error_u_vector4[59] + error_u_vector4[60] + error_u_vector4[61] + error_u_vector4[62] + error_u_vector4[63] + error_u_vector4[64] + error_u_vector4[65] + error_u_vector4[66] + error_u_vector4[67] + error_u_vector4[68] + error_u_vector4[69] + error_u_vector4[70] + error_u_vector4[71] + error_u_vector4[72] + error_u_vector4[73] + error_u_vector4[74] + error_u_vector4[75] + error_u_vector4[76] + error_u_vector4[77] + error_u_vector4[78] + error_u_vector4[79] + error_u_vector4[80] + error_u_vector4[81] + error_u_vector4[82] + error_u_vector4[83] + error_u_vector4[84] + error_u_vector4[85] + error_u_vector4[86] + error_u_vector4[87] + error_u_vector4[88] + error_u_vector4[89] + error_u_vector4[90] + error_u_vector4[91] + error_u_vector4[92] + error_u_vector4[93] + error_u_vector4[94] + error_u_vector4[95] + error_u_vector4[96] + error_u_vector4[97] + error_u_vector4[98] + error_u_vector4[99] + error_u_vector4[100] + error_u_vector4[101] + error_u_vector4[102] + error_u_vector4[103] + error_u_vector4[104] + error_u_vector4[105] + error_u_vector4[106] + error_u_vector4[107] + error_u_vector4[108] + error_u_vector4[109] + error_u_vector4[110] + error_u_vector4[111] + error_u_vector4[112] + error_u_vector4[113] + error_u_vector4[114] + error_u_vector4[115] + error_u_vector4[116] + error_u_vector4[117] + error_u_vector4[118] + error_u_vector4[119] + error_u_vector4[120] + error_u_vector4[121] + error_u_vector4[122] + error_u_vector4[123] + error_u_vector4[124] + error_u_vector4[125] + error_u_vector4[126] + error_u_vector4[127] + error_u_vector4[128] + error_u_vector4[129] + error_u_vector4[130] + error_u_vector4[131] + error_u_vector4[132] + error_u_vector4[133] + error_u_vector4[134] + error_u_vector4[135] + error_u_vector4[136] + error_u_vector4[137] + error_u_vector4[138] + error_u_vector4[139] + error_u_vector4[140] + error_u_vector4[141] + error_u_vector4[142] + error_u_vector4[143] + error_u_vector4[144] + error_u_vector4[145] + error_u_vector4[146] + error_u_vector4[147] + error_u_vector4[148] + error_u_vector4[149] + error_u_vector4[150] + error_u_vector4[151] + error_u_vector4[152] + error_u_vector4[153] + error_u_vector4[154] + error_u_vector4[155] + error_u_vector4[156] + error_u_vector4[157] + error_u_vector4[158] + error_u_vector4[159] + error_u_vector4[160] + error_u_vector4[161] + error_u_vector4[162] + error_u_vector4[163] + error_u_vector4[164] + error_u_vector4[165] + error_u_vector4[166] + error_u_vector4[167] + error_u_vector4[168] + error_u_vector4[169] + error_u_vector4[170] + error_u_vector4[171] + error_u_vector4[172] + error_u_vector4[173] + error_u_vector4[174] + error_u_vector4[175] + error_u_vector4[176] + error_u_vector4[177] + error_u_vector4[178] + error_u_vector4[179] + error_u_vector4[180] + error_u_vector4[181] + error_u_vector4[182] + error_u_vector4[183] + error_u_vector4[184] + error_u_vector4[185] + error_u_vector4[186] + error_u_vector4[187] + error_u_vector4[188] + error_u_vector4[189] + error_u_vector4[190] + error_u_vector4[191] + error_u_vector4[192] + error_u_vector4[193] + error_u_vector4[194] + error_u_vector4[195] + error_u_vector4[196] + error_u_vector4[197] + error_u_vector4[198] + error_u_vector4[199] + error_u_vector4[200] + error_u_vector4[201] + error_u_vector4[202] + error_u_vector4[203] + error_u_vector4[204] + error_u_vector4[205] + error_u_vector4[206] + error_u_vector4[207] + error_u_vector4[208] + error_u_vector4[209] + error_u_vector4[210] + error_u_vector4[211] + error_u_vector4[212] + error_u_vector4[213] + error_u_vector4[214] + error_u_vector4[215] + error_u_vector4[216] + error_u_vector4[217] + error_u_vector4[218] + error_u_vector4[219] + error_u_vector4[220] + error_u_vector4[221] + error_u_vector4[222] + error_u_vector4[223] + error_u_vector4[224] + error_u_vector4[225] + error_u_vector4[226] + error_u_vector4[227] + error_u_vector4[228] + error_u_vector4[229] + error_u_vector4[230] + error_u_vector4[231] + error_u_vector4[232] + error_u_vector4[233] + error_u_vector4[234] + error_u_vector4[235] + error_u_vector4[236] + error_u_vector4[237] + error_u_vector4[238]; 
            errs5_u <= error_u_vector5[0] + error_u_vector5[1] + error_u_vector5[2] + error_u_vector5[3] + error_u_vector5[4] + error_u_vector5[5] + error_u_vector5[6] + error_u_vector5[7] + error_u_vector5[8] + error_u_vector5[9] + error_u_vector5[10] + error_u_vector5[11] + error_u_vector5[12] + error_u_vector5[13] + error_u_vector5[14] + error_u_vector5[15] + error_u_vector5[16] + error_u_vector5[17] + error_u_vector5[18] + error_u_vector5[19] + error_u_vector5[20] + error_u_vector5[21] + error_u_vector5[22] + error_u_vector5[23] + error_u_vector5[24] + error_u_vector5[25] + error_u_vector5[26] + error_u_vector5[27] + error_u_vector5[28] + error_u_vector5[29] + error_u_vector5[30] + error_u_vector5[31] + error_u_vector5[32] + error_u_vector5[33] + error_u_vector5[34] + error_u_vector5[35] + error_u_vector5[36] + error_u_vector5[37] + error_u_vector5[38] + error_u_vector5[39] + error_u_vector5[40] + error_u_vector5[41] + error_u_vector5[42] + error_u_vector5[43] + error_u_vector5[44] + error_u_vector5[45] + error_u_vector5[46] + error_u_vector5[47] + error_u_vector5[48] + error_u_vector5[49] + error_u_vector5[50] + error_u_vector5[51] + error_u_vector5[52] + error_u_vector5[53] + error_u_vector5[54] + error_u_vector5[55] + error_u_vector5[56] + error_u_vector5[57] + error_u_vector5[58] + error_u_vector5[59] + error_u_vector5[60] + error_u_vector5[61] + error_u_vector5[62] + error_u_vector5[63] + error_u_vector5[64] + error_u_vector5[65] + error_u_vector5[66] + error_u_vector5[67] + error_u_vector5[68] + error_u_vector5[69] + error_u_vector5[70] + error_u_vector5[71] + error_u_vector5[72] + error_u_vector5[73] + error_u_vector5[74] + error_u_vector5[75] + error_u_vector5[76] + error_u_vector5[77] + error_u_vector5[78] + error_u_vector5[79] + error_u_vector5[80] + error_u_vector5[81] + error_u_vector5[82] + error_u_vector5[83] + error_u_vector5[84] + error_u_vector5[85] + error_u_vector5[86] + error_u_vector5[87] + error_u_vector5[88] + error_u_vector5[89] + error_u_vector5[90] + error_u_vector5[91] + error_u_vector5[92] + error_u_vector5[93] + error_u_vector5[94] + error_u_vector5[95] + error_u_vector5[96] + error_u_vector5[97] + error_u_vector5[98] + error_u_vector5[99] + error_u_vector5[100] + error_u_vector5[101] + error_u_vector5[102] + error_u_vector5[103] + error_u_vector5[104] + error_u_vector5[105] + error_u_vector5[106] + error_u_vector5[107] + error_u_vector5[108] + error_u_vector5[109] + error_u_vector5[110] + error_u_vector5[111] + error_u_vector5[112] + error_u_vector5[113] + error_u_vector5[114] + error_u_vector5[115] + error_u_vector5[116] + error_u_vector5[117] + error_u_vector5[118] + error_u_vector5[119] + error_u_vector5[120] + error_u_vector5[121] + error_u_vector5[122] + error_u_vector5[123] + error_u_vector5[124] + error_u_vector5[125] + error_u_vector5[126] + error_u_vector5[127] + error_u_vector5[128] + error_u_vector5[129] + error_u_vector5[130] + error_u_vector5[131] + error_u_vector5[132] + error_u_vector5[133] + error_u_vector5[134] + error_u_vector5[135] + error_u_vector5[136] + error_u_vector5[137] + error_u_vector5[138] + error_u_vector5[139] + error_u_vector5[140] + error_u_vector5[141] + error_u_vector5[142] + error_u_vector5[143] + error_u_vector5[144] + error_u_vector5[145] + error_u_vector5[146] + error_u_vector5[147] + error_u_vector5[148] + error_u_vector5[149] + error_u_vector5[150] + error_u_vector5[151] + error_u_vector5[152] + error_u_vector5[153] + error_u_vector5[154] + error_u_vector5[155] + error_u_vector5[156] + error_u_vector5[157] + error_u_vector5[158] + error_u_vector5[159] + error_u_vector5[160] + error_u_vector5[161] + error_u_vector5[162] + error_u_vector5[163] + error_u_vector5[164] + error_u_vector5[165] + error_u_vector5[166] + error_u_vector5[167] + error_u_vector5[168] + error_u_vector5[169] + error_u_vector5[170] + error_u_vector5[171] + error_u_vector5[172] + error_u_vector5[173] + error_u_vector5[174] + error_u_vector5[175] + error_u_vector5[176] + error_u_vector5[177] + error_u_vector5[178] + error_u_vector5[179] + error_u_vector5[180] + error_u_vector5[181] + error_u_vector5[182] + error_u_vector5[183] + error_u_vector5[184] + error_u_vector5[185] + error_u_vector5[186] + error_u_vector5[187] + error_u_vector5[188] + error_u_vector5[189] + error_u_vector5[190] + error_u_vector5[191] + error_u_vector5[192] + error_u_vector5[193] + error_u_vector5[194] + error_u_vector5[195] + error_u_vector5[196] + error_u_vector5[197] + error_u_vector5[198] + error_u_vector5[199] + error_u_vector5[200] + error_u_vector5[201] + error_u_vector5[202] + error_u_vector5[203] + error_u_vector5[204] + error_u_vector5[205] + error_u_vector5[206] + error_u_vector5[207] + error_u_vector5[208] + error_u_vector5[209] + error_u_vector5[210] + error_u_vector5[211] + error_u_vector5[212] + error_u_vector5[213] + error_u_vector5[214] + error_u_vector5[215] + error_u_vector5[216] + error_u_vector5[217] + error_u_vector5[218] + error_u_vector5[219] + error_u_vector5[220] + error_u_vector5[221] + error_u_vector5[222] + error_u_vector5[223] + error_u_vector5[224] + error_u_vector5[225] + error_u_vector5[226] + error_u_vector5[227] + error_u_vector5[228] + error_u_vector5[229] + error_u_vector5[230] + error_u_vector5[231] + error_u_vector5[232] + error_u_vector5[233] + error_u_vector5[234] + error_u_vector5[235] + error_u_vector5[236] + error_u_vector5[237] + error_u_vector5[238]; 
            errs6_u <= error_u_vector6[0] + error_u_vector6[1] + error_u_vector6[2] + error_u_vector6[3] + error_u_vector6[4] + error_u_vector6[5] + error_u_vector6[6] + error_u_vector6[7] + error_u_vector6[8] + error_u_vector6[9] + error_u_vector6[10] + error_u_vector6[11] + error_u_vector6[12] + error_u_vector6[13] + error_u_vector6[14] + error_u_vector6[15] + error_u_vector6[16] + error_u_vector6[17] + error_u_vector6[18] + error_u_vector6[19] + error_u_vector6[20] + error_u_vector6[21] + error_u_vector6[22] + error_u_vector6[23] + error_u_vector6[24] + error_u_vector6[25] + error_u_vector6[26] + error_u_vector6[27] + error_u_vector6[28] + error_u_vector6[29] + error_u_vector6[30] + error_u_vector6[31] + error_u_vector6[32] + error_u_vector6[33] + error_u_vector6[34] + error_u_vector6[35] + error_u_vector6[36] + error_u_vector6[37] + error_u_vector6[38] + error_u_vector6[39] + error_u_vector6[40] + error_u_vector6[41] + error_u_vector6[42] + error_u_vector6[43] + error_u_vector6[44] + error_u_vector6[45] + error_u_vector6[46] + error_u_vector6[47] + error_u_vector6[48] + error_u_vector6[49] + error_u_vector6[50] + error_u_vector6[51] + error_u_vector6[52] + error_u_vector6[53] + error_u_vector6[54] + error_u_vector6[55] + error_u_vector6[56] + error_u_vector6[57] + error_u_vector6[58] + error_u_vector6[59] + error_u_vector6[60] + error_u_vector6[61] + error_u_vector6[62] + error_u_vector6[63] + error_u_vector6[64] + error_u_vector6[65] + error_u_vector6[66] + error_u_vector6[67] + error_u_vector6[68] + error_u_vector6[69] + error_u_vector6[70] + error_u_vector6[71] + error_u_vector6[72] + error_u_vector6[73] + error_u_vector6[74] + error_u_vector6[75] + error_u_vector6[76] + error_u_vector6[77] + error_u_vector6[78] + error_u_vector6[79] + error_u_vector6[80] + error_u_vector6[81] + error_u_vector6[82] + error_u_vector6[83] + error_u_vector6[84] + error_u_vector6[85] + error_u_vector6[86] + error_u_vector6[87] + error_u_vector6[88] + error_u_vector6[89] + error_u_vector6[90] + error_u_vector6[91] + error_u_vector6[92] + error_u_vector6[93] + error_u_vector6[94] + error_u_vector6[95] + error_u_vector6[96] + error_u_vector6[97] + error_u_vector6[98] + error_u_vector6[99] + error_u_vector6[100] + error_u_vector6[101] + error_u_vector6[102] + error_u_vector6[103] + error_u_vector6[104] + error_u_vector6[105] + error_u_vector6[106] + error_u_vector6[107] + error_u_vector6[108] + error_u_vector6[109] + error_u_vector6[110] + error_u_vector6[111] + error_u_vector6[112] + error_u_vector6[113] + error_u_vector6[114] + error_u_vector6[115] + error_u_vector6[116] + error_u_vector6[117] + error_u_vector6[118] + error_u_vector6[119] + error_u_vector6[120] + error_u_vector6[121] + error_u_vector6[122] + error_u_vector6[123] + error_u_vector6[124] + error_u_vector6[125] + error_u_vector6[126] + error_u_vector6[127] + error_u_vector6[128] + error_u_vector6[129] + error_u_vector6[130] + error_u_vector6[131] + error_u_vector6[132] + error_u_vector6[133] + error_u_vector6[134] + error_u_vector6[135] + error_u_vector6[136] + error_u_vector6[137] + error_u_vector6[138] + error_u_vector6[139] + error_u_vector6[140] + error_u_vector6[141] + error_u_vector6[142] + error_u_vector6[143] + error_u_vector6[144] + error_u_vector6[145] + error_u_vector6[146] + error_u_vector6[147] + error_u_vector6[148] + error_u_vector6[149] + error_u_vector6[150] + error_u_vector6[151] + error_u_vector6[152] + error_u_vector6[153] + error_u_vector6[154] + error_u_vector6[155] + error_u_vector6[156] + error_u_vector6[157] + error_u_vector6[158] + error_u_vector6[159] + error_u_vector6[160] + error_u_vector6[161] + error_u_vector6[162] + error_u_vector6[163] + error_u_vector6[164] + error_u_vector6[165] + error_u_vector6[166] + error_u_vector6[167] + error_u_vector6[168] + error_u_vector6[169] + error_u_vector6[170] + error_u_vector6[171] + error_u_vector6[172] + error_u_vector6[173] + error_u_vector6[174] + error_u_vector6[175] + error_u_vector6[176] + error_u_vector6[177] + error_u_vector6[178] + error_u_vector6[179] + error_u_vector6[180] + error_u_vector6[181] + error_u_vector6[182] + error_u_vector6[183] + error_u_vector6[184] + error_u_vector6[185] + error_u_vector6[186] + error_u_vector6[187] + error_u_vector6[188] + error_u_vector6[189] + error_u_vector6[190] + error_u_vector6[191] + error_u_vector6[192] + error_u_vector6[193] + error_u_vector6[194] + error_u_vector6[195] + error_u_vector6[196] + error_u_vector6[197] + error_u_vector6[198] + error_u_vector6[199] + error_u_vector6[200] + error_u_vector6[201] + error_u_vector6[202] + error_u_vector6[203] + error_u_vector6[204] + error_u_vector6[205] + error_u_vector6[206] + error_u_vector6[207] + error_u_vector6[208] + error_u_vector6[209] + error_u_vector6[210] + error_u_vector6[211] + error_u_vector6[212] + error_u_vector6[213] + error_u_vector6[214] + error_u_vector6[215] + error_u_vector6[216] + error_u_vector6[217] + error_u_vector6[218] + error_u_vector6[219] + error_u_vector6[220] + error_u_vector6[221] + error_u_vector6[222] + error_u_vector6[223] + error_u_vector6[224] + error_u_vector6[225] + error_u_vector6[226] + error_u_vector6[227] + error_u_vector6[228] + error_u_vector6[229] + error_u_vector6[230] + error_u_vector6[231] + error_u_vector6[232] + error_u_vector6[233] + error_u_vector6[234] + error_u_vector6[235] + error_u_vector6[236] + error_u_vector6[237] + error_u_vector6[238]; 
            errs7_u <= error_u_vector7[0] + error_u_vector7[1] + error_u_vector7[2] + error_u_vector7[3] + error_u_vector7[4] + error_u_vector7[5] + error_u_vector7[6] + error_u_vector7[7] + error_u_vector7[8] + error_u_vector7[9] + error_u_vector7[10] + error_u_vector7[11] + error_u_vector7[12] + error_u_vector7[13] + error_u_vector7[14] + error_u_vector7[15] + error_u_vector7[16] + error_u_vector7[17] + error_u_vector7[18] + error_u_vector7[19] + error_u_vector7[20] + error_u_vector7[21] + error_u_vector7[22] + error_u_vector7[23] + error_u_vector7[24] + error_u_vector7[25] + error_u_vector7[26] + error_u_vector7[27] + error_u_vector7[28] + error_u_vector7[29] + error_u_vector7[30] + error_u_vector7[31] + error_u_vector7[32] + error_u_vector7[33] + error_u_vector7[34] + error_u_vector7[35] + error_u_vector7[36] + error_u_vector7[37] + error_u_vector7[38] + error_u_vector7[39] + error_u_vector7[40] + error_u_vector7[41] + error_u_vector7[42] + error_u_vector7[43] + error_u_vector7[44] + error_u_vector7[45] + error_u_vector7[46] + error_u_vector7[47] + error_u_vector7[48] + error_u_vector7[49] + error_u_vector7[50] + error_u_vector7[51] + error_u_vector7[52] + error_u_vector7[53] + error_u_vector7[54] + error_u_vector7[55] + error_u_vector7[56] + error_u_vector7[57] + error_u_vector7[58] + error_u_vector7[59] + error_u_vector7[60] + error_u_vector7[61] + error_u_vector7[62] + error_u_vector7[63] + error_u_vector7[64] + error_u_vector7[65] + error_u_vector7[66] + error_u_vector7[67] + error_u_vector7[68] + error_u_vector7[69] + error_u_vector7[70] + error_u_vector7[71] + error_u_vector7[72] + error_u_vector7[73] + error_u_vector7[74] + error_u_vector7[75] + error_u_vector7[76] + error_u_vector7[77] + error_u_vector7[78] + error_u_vector7[79] + error_u_vector7[80] + error_u_vector7[81] + error_u_vector7[82] + error_u_vector7[83] + error_u_vector7[84] + error_u_vector7[85] + error_u_vector7[86] + error_u_vector7[87] + error_u_vector7[88] + error_u_vector7[89] + error_u_vector7[90] + error_u_vector7[91] + error_u_vector7[92] + error_u_vector7[93] + error_u_vector7[94] + error_u_vector7[95] + error_u_vector7[96] + error_u_vector7[97] + error_u_vector7[98] + error_u_vector7[99] + error_u_vector7[100] + error_u_vector7[101] + error_u_vector7[102] + error_u_vector7[103] + error_u_vector7[104] + error_u_vector7[105] + error_u_vector7[106] + error_u_vector7[107] + error_u_vector7[108] + error_u_vector7[109] + error_u_vector7[110] + error_u_vector7[111] + error_u_vector7[112] + error_u_vector7[113] + error_u_vector7[114] + error_u_vector7[115] + error_u_vector7[116] + error_u_vector7[117] + error_u_vector7[118] + error_u_vector7[119] + error_u_vector7[120] + error_u_vector7[121] + error_u_vector7[122] + error_u_vector7[123] + error_u_vector7[124] + error_u_vector7[125] + error_u_vector7[126] + error_u_vector7[127] + error_u_vector7[128] + error_u_vector7[129] + error_u_vector7[130] + error_u_vector7[131] + error_u_vector7[132] + error_u_vector7[133] + error_u_vector7[134] + error_u_vector7[135] + error_u_vector7[136] + error_u_vector7[137] + error_u_vector7[138] + error_u_vector7[139] + error_u_vector7[140] + error_u_vector7[141] + error_u_vector7[142] + error_u_vector7[143] + error_u_vector7[144] + error_u_vector7[145] + error_u_vector7[146] + error_u_vector7[147] + error_u_vector7[148] + error_u_vector7[149] + error_u_vector7[150] + error_u_vector7[151] + error_u_vector7[152] + error_u_vector7[153] + error_u_vector7[154] + error_u_vector7[155] + error_u_vector7[156] + error_u_vector7[157] + error_u_vector7[158] + error_u_vector7[159] + error_u_vector7[160] + error_u_vector7[161] + error_u_vector7[162] + error_u_vector7[163] + error_u_vector7[164] + error_u_vector7[165] + error_u_vector7[166] + error_u_vector7[167] + error_u_vector7[168] + error_u_vector7[169] + error_u_vector7[170] + error_u_vector7[171] + error_u_vector7[172] + error_u_vector7[173] + error_u_vector7[174] + error_u_vector7[175] + error_u_vector7[176] + error_u_vector7[177] + error_u_vector7[178] + error_u_vector7[179] + error_u_vector7[180] + error_u_vector7[181] + error_u_vector7[182] + error_u_vector7[183] + error_u_vector7[184] + error_u_vector7[185] + error_u_vector7[186] + error_u_vector7[187] + error_u_vector7[188] + error_u_vector7[189] + error_u_vector7[190] + error_u_vector7[191] + error_u_vector7[192] + error_u_vector7[193] + error_u_vector7[194] + error_u_vector7[195] + error_u_vector7[196] + error_u_vector7[197] + error_u_vector7[198] + error_u_vector7[199] + error_u_vector7[200] + error_u_vector7[201] + error_u_vector7[202] + error_u_vector7[203] + error_u_vector7[204] + error_u_vector7[205] + error_u_vector7[206] + error_u_vector7[207] + error_u_vector7[208] + error_u_vector7[209] + error_u_vector7[210] + error_u_vector7[211] + error_u_vector7[212] + error_u_vector7[213] + error_u_vector7[214] + error_u_vector7[215] + error_u_vector7[216] + error_u_vector7[217] + error_u_vector7[218] + error_u_vector7[219] + error_u_vector7[220] + error_u_vector7[221] + error_u_vector7[222] + error_u_vector7[223] + error_u_vector7[224] + error_u_vector7[225] + error_u_vector7[226] + error_u_vector7[227] + error_u_vector7[228] + error_u_vector7[229] + error_u_vector7[230] + error_u_vector7[231] + error_u_vector7[232] + error_u_vector7[233] + error_u_vector7[234] + error_u_vector7[235] + error_u_vector7[236] + error_u_vector7[237] + error_u_vector7[238]; 
            errs8_u <= error_u_vector8[0] + error_u_vector8[1] + error_u_vector8[2] + error_u_vector8[3] + error_u_vector8[4] + error_u_vector8[5] + error_u_vector8[6] + error_u_vector8[7] + error_u_vector8[8] + error_u_vector8[9] + error_u_vector8[10] + error_u_vector8[11] + error_u_vector8[12] + error_u_vector8[13] + error_u_vector8[14] + error_u_vector8[15] + error_u_vector8[16] + error_u_vector8[17] + error_u_vector8[18] + error_u_vector8[19] + error_u_vector8[20] + error_u_vector8[21] + error_u_vector8[22] + error_u_vector8[23] + error_u_vector8[24] + error_u_vector8[25] + error_u_vector8[26] + error_u_vector8[27] + error_u_vector8[28] + error_u_vector8[29] + error_u_vector8[30] + error_u_vector8[31] + error_u_vector8[32] + error_u_vector8[33] + error_u_vector8[34] + error_u_vector8[35] + error_u_vector8[36] + error_u_vector8[37] + error_u_vector8[38] + error_u_vector8[39] + error_u_vector8[40] + error_u_vector8[41] + error_u_vector8[42] + error_u_vector8[43] + error_u_vector8[44] + error_u_vector8[45] + error_u_vector8[46] + error_u_vector8[47] + error_u_vector8[48] + error_u_vector8[49] + error_u_vector8[50] + error_u_vector8[51] + error_u_vector8[52] + error_u_vector8[53] + error_u_vector8[54] + error_u_vector8[55] + error_u_vector8[56] + error_u_vector8[57] + error_u_vector8[58] + error_u_vector8[59] + error_u_vector8[60] + error_u_vector8[61] + error_u_vector8[62] + error_u_vector8[63] + error_u_vector8[64] + error_u_vector8[65] + error_u_vector8[66] + error_u_vector8[67] + error_u_vector8[68] + error_u_vector8[69] + error_u_vector8[70] + error_u_vector8[71] + error_u_vector8[72] + error_u_vector8[73] + error_u_vector8[74] + error_u_vector8[75] + error_u_vector8[76] + error_u_vector8[77] + error_u_vector8[78] + error_u_vector8[79] + error_u_vector8[80] + error_u_vector8[81] + error_u_vector8[82] + error_u_vector8[83] + error_u_vector8[84] + error_u_vector8[85] + error_u_vector8[86] + error_u_vector8[87] + error_u_vector8[88] + error_u_vector8[89] + error_u_vector8[90] + error_u_vector8[91] + error_u_vector8[92] + error_u_vector8[93] + error_u_vector8[94] + error_u_vector8[95] + error_u_vector8[96] + error_u_vector8[97] + error_u_vector8[98] + error_u_vector8[99] + error_u_vector8[100] + error_u_vector8[101] + error_u_vector8[102] + error_u_vector8[103] + error_u_vector8[104] + error_u_vector8[105] + error_u_vector8[106] + error_u_vector8[107] + error_u_vector8[108] + error_u_vector8[109] + error_u_vector8[110] + error_u_vector8[111] + error_u_vector8[112] + error_u_vector8[113] + error_u_vector8[114] + error_u_vector8[115] + error_u_vector8[116] + error_u_vector8[117] + error_u_vector8[118] + error_u_vector8[119] + error_u_vector8[120] + error_u_vector8[121] + error_u_vector8[122] + error_u_vector8[123] + error_u_vector8[124] + error_u_vector8[125] + error_u_vector8[126] + error_u_vector8[127] + error_u_vector8[128] + error_u_vector8[129] + error_u_vector8[130] + error_u_vector8[131] + error_u_vector8[132] + error_u_vector8[133] + error_u_vector8[134] + error_u_vector8[135] + error_u_vector8[136] + error_u_vector8[137] + error_u_vector8[138] + error_u_vector8[139] + error_u_vector8[140] + error_u_vector8[141] + error_u_vector8[142] + error_u_vector8[143] + error_u_vector8[144] + error_u_vector8[145] + error_u_vector8[146] + error_u_vector8[147] + error_u_vector8[148] + error_u_vector8[149] + error_u_vector8[150] + error_u_vector8[151] + error_u_vector8[152] + error_u_vector8[153] + error_u_vector8[154] + error_u_vector8[155] + error_u_vector8[156] + error_u_vector8[157] + error_u_vector8[158] + error_u_vector8[159] + error_u_vector8[160] + error_u_vector8[161] + error_u_vector8[162] + error_u_vector8[163] + error_u_vector8[164] + error_u_vector8[165] + error_u_vector8[166] + error_u_vector8[167] + error_u_vector8[168] + error_u_vector8[169] + error_u_vector8[170] + error_u_vector8[171] + error_u_vector8[172] + error_u_vector8[173] + error_u_vector8[174] + error_u_vector8[175] + error_u_vector8[176] + error_u_vector8[177] + error_u_vector8[178] + error_u_vector8[179] + error_u_vector8[180] + error_u_vector8[181] + error_u_vector8[182] + error_u_vector8[183] + error_u_vector8[184] + error_u_vector8[185] + error_u_vector8[186] + error_u_vector8[187] + error_u_vector8[188] + error_u_vector8[189] + error_u_vector8[190] + error_u_vector8[191] + error_u_vector8[192] + error_u_vector8[193] + error_u_vector8[194] + error_u_vector8[195] + error_u_vector8[196] + error_u_vector8[197] + error_u_vector8[198] + error_u_vector8[199] + error_u_vector8[200] + error_u_vector8[201] + error_u_vector8[202] + error_u_vector8[203] + error_u_vector8[204] + error_u_vector8[205] + error_u_vector8[206] + error_u_vector8[207] + error_u_vector8[208] + error_u_vector8[209] + error_u_vector8[210] + error_u_vector8[211] + error_u_vector8[212] + error_u_vector8[213] + error_u_vector8[214] + error_u_vector8[215] + error_u_vector8[216] + error_u_vector8[217] + error_u_vector8[218] + error_u_vector8[219] + error_u_vector8[220] + error_u_vector8[221] + error_u_vector8[222] + error_u_vector8[223] + error_u_vector8[224] + error_u_vector8[225] + error_u_vector8[226] + error_u_vector8[227] + error_u_vector8[228] + error_u_vector8[229] + error_u_vector8[230] + error_u_vector8[231] + error_u_vector8[232] + error_u_vector8[233] + error_u_vector8[234] + error_u_vector8[235] + error_u_vector8[236] + error_u_vector8[237] + error_u_vector8[238]; 
            errs9_u <= error_u_vector9[0] + error_u_vector9[1] + error_u_vector9[2] + error_u_vector9[3] + error_u_vector9[4] + error_u_vector9[5] + error_u_vector9[6] + error_u_vector9[7] + error_u_vector9[8] + error_u_vector9[9] + error_u_vector9[10] + error_u_vector9[11] + error_u_vector9[12] + error_u_vector9[13] + error_u_vector9[14] + error_u_vector9[15] + error_u_vector9[16] + error_u_vector9[17] + error_u_vector9[18] + error_u_vector9[19] + error_u_vector9[20] + error_u_vector9[21] + error_u_vector9[22] + error_u_vector9[23] + error_u_vector9[24] + error_u_vector9[25] + error_u_vector9[26] + error_u_vector9[27] + error_u_vector9[28] + error_u_vector9[29] + error_u_vector9[30] + error_u_vector9[31] + error_u_vector9[32] + error_u_vector9[33] + error_u_vector9[34] + error_u_vector9[35] + error_u_vector9[36] + error_u_vector9[37] + error_u_vector9[38] + error_u_vector9[39] + error_u_vector9[40] + error_u_vector9[41] + error_u_vector9[42] + error_u_vector9[43] + error_u_vector9[44] + error_u_vector9[45] + error_u_vector9[46] + error_u_vector9[47] + error_u_vector9[48] + error_u_vector9[49] + error_u_vector9[50] + error_u_vector9[51] + error_u_vector9[52] + error_u_vector9[53] + error_u_vector9[54] + error_u_vector9[55] + error_u_vector9[56] + error_u_vector9[57] + error_u_vector9[58] + error_u_vector9[59] + error_u_vector9[60] + error_u_vector9[61] + error_u_vector9[62] + error_u_vector9[63] + error_u_vector9[64] + error_u_vector9[65] + error_u_vector9[66] + error_u_vector9[67] + error_u_vector9[68] + error_u_vector9[69] + error_u_vector9[70] + error_u_vector9[71] + error_u_vector9[72] + error_u_vector9[73] + error_u_vector9[74] + error_u_vector9[75] + error_u_vector9[76] + error_u_vector9[77] + error_u_vector9[78] + error_u_vector9[79] + error_u_vector9[80] + error_u_vector9[81] + error_u_vector9[82] + error_u_vector9[83] + error_u_vector9[84] + error_u_vector9[85] + error_u_vector9[86] + error_u_vector9[87] + error_u_vector9[88] + error_u_vector9[89] + error_u_vector9[90] + error_u_vector9[91] + error_u_vector9[92] + error_u_vector9[93] + error_u_vector9[94] + error_u_vector9[95] + error_u_vector9[96] + error_u_vector9[97] + error_u_vector9[98] + error_u_vector9[99] + error_u_vector9[100] + error_u_vector9[101] + error_u_vector9[102] + error_u_vector9[103] + error_u_vector9[104] + error_u_vector9[105] + error_u_vector9[106] + error_u_vector9[107] + error_u_vector9[108] + error_u_vector9[109] + error_u_vector9[110] + error_u_vector9[111] + error_u_vector9[112] + error_u_vector9[113] + error_u_vector9[114] + error_u_vector9[115] + error_u_vector9[116] + error_u_vector9[117] + error_u_vector9[118] + error_u_vector9[119] + error_u_vector9[120] + error_u_vector9[121] + error_u_vector9[122] + error_u_vector9[123] + error_u_vector9[124] + error_u_vector9[125] + error_u_vector9[126] + error_u_vector9[127] + error_u_vector9[128] + error_u_vector9[129] + error_u_vector9[130] + error_u_vector9[131] + error_u_vector9[132] + error_u_vector9[133] + error_u_vector9[134] + error_u_vector9[135] + error_u_vector9[136] + error_u_vector9[137] + error_u_vector9[138] + error_u_vector9[139] + error_u_vector9[140] + error_u_vector9[141] + error_u_vector9[142] + error_u_vector9[143] + error_u_vector9[144] + error_u_vector9[145] + error_u_vector9[146] + error_u_vector9[147] + error_u_vector9[148] + error_u_vector9[149] + error_u_vector9[150] + error_u_vector9[151] + error_u_vector9[152] + error_u_vector9[153] + error_u_vector9[154] + error_u_vector9[155] + error_u_vector9[156] + error_u_vector9[157] + error_u_vector9[158] + error_u_vector9[159] + error_u_vector9[160] + error_u_vector9[161] + error_u_vector9[162] + error_u_vector9[163] + error_u_vector9[164] + error_u_vector9[165] + error_u_vector9[166] + error_u_vector9[167] + error_u_vector9[168] + error_u_vector9[169] + error_u_vector9[170] + error_u_vector9[171] + error_u_vector9[172] + error_u_vector9[173] + error_u_vector9[174] + error_u_vector9[175] + error_u_vector9[176] + error_u_vector9[177] + error_u_vector9[178] + error_u_vector9[179] + error_u_vector9[180] + error_u_vector9[181] + error_u_vector9[182] + error_u_vector9[183] + error_u_vector9[184] + error_u_vector9[185] + error_u_vector9[186] + error_u_vector9[187] + error_u_vector9[188] + error_u_vector9[189] + error_u_vector9[190] + error_u_vector9[191] + error_u_vector9[192] + error_u_vector9[193] + error_u_vector9[194] + error_u_vector9[195] + error_u_vector9[196] + error_u_vector9[197] + error_u_vector9[198] + error_u_vector9[199] + error_u_vector9[200] + error_u_vector9[201] + error_u_vector9[202] + error_u_vector9[203] + error_u_vector9[204] + error_u_vector9[205] + error_u_vector9[206] + error_u_vector9[207] + error_u_vector9[208] + error_u_vector9[209] + error_u_vector9[210] + error_u_vector9[211] + error_u_vector9[212] + error_u_vector9[213] + error_u_vector9[214] + error_u_vector9[215] + error_u_vector9[216] + error_u_vector9[217] + error_u_vector9[218] + error_u_vector9[219] + error_u_vector9[220] + error_u_vector9[221] + error_u_vector9[222] + error_u_vector9[223] + error_u_vector9[224] + error_u_vector9[225] + error_u_vector9[226] + error_u_vector9[227] + error_u_vector9[228] + error_u_vector9[229] + error_u_vector9[230] + error_u_vector9[231] + error_u_vector9[232] + error_u_vector9[233] + error_u_vector9[234] + error_u_vector9[235] + error_u_vector9[236] + error_u_vector9[237] + error_u_vector9[238]; 
            errs10_u <= error_u_vector10[0] + error_u_vector10[1] + error_u_vector10[2] + error_u_vector10[3] + error_u_vector10[4] + error_u_vector10[5] + error_u_vector10[6] + error_u_vector10[7] + error_u_vector10[8] + error_u_vector10[9] + error_u_vector10[10] + error_u_vector10[11] + error_u_vector10[12] + error_u_vector10[13] + error_u_vector10[14] + error_u_vector10[15] + error_u_vector10[16] + error_u_vector10[17] + error_u_vector10[18] + error_u_vector10[19] + error_u_vector10[20] + error_u_vector10[21] + error_u_vector10[22] + error_u_vector10[23] + error_u_vector10[24] + error_u_vector10[25] + error_u_vector10[26] + error_u_vector10[27] + error_u_vector10[28] + error_u_vector10[29] + error_u_vector10[30] + error_u_vector10[31] + error_u_vector10[32] + error_u_vector10[33] + error_u_vector10[34] + error_u_vector10[35] + error_u_vector10[36] + error_u_vector10[37] + error_u_vector10[38] + error_u_vector10[39] + error_u_vector10[40] + error_u_vector10[41] + error_u_vector10[42] + error_u_vector10[43] + error_u_vector10[44] + error_u_vector10[45] + error_u_vector10[46] + error_u_vector10[47] + error_u_vector10[48] + error_u_vector10[49] + error_u_vector10[50] + error_u_vector10[51] + error_u_vector10[52] + error_u_vector10[53] + error_u_vector10[54] + error_u_vector10[55] + error_u_vector10[56] + error_u_vector10[57] + error_u_vector10[58] + error_u_vector10[59] + error_u_vector10[60] + error_u_vector10[61] + error_u_vector10[62] + error_u_vector10[63] + error_u_vector10[64] + error_u_vector10[65] + error_u_vector10[66] + error_u_vector10[67] + error_u_vector10[68] + error_u_vector10[69] + error_u_vector10[70] + error_u_vector10[71] + error_u_vector10[72] + error_u_vector10[73] + error_u_vector10[74] + error_u_vector10[75] + error_u_vector10[76] + error_u_vector10[77] + error_u_vector10[78] + error_u_vector10[79] + error_u_vector10[80] + error_u_vector10[81] + error_u_vector10[82] + error_u_vector10[83] + error_u_vector10[84] + error_u_vector10[85] + error_u_vector10[86] + error_u_vector10[87] + error_u_vector10[88] + error_u_vector10[89] + error_u_vector10[90] + error_u_vector10[91] + error_u_vector10[92] + error_u_vector10[93] + error_u_vector10[94] + error_u_vector10[95] + error_u_vector10[96] + error_u_vector10[97] + error_u_vector10[98] + error_u_vector10[99] + error_u_vector10[100] + error_u_vector10[101] + error_u_vector10[102] + error_u_vector10[103] + error_u_vector10[104] + error_u_vector10[105] + error_u_vector10[106] + error_u_vector10[107] + error_u_vector10[108] + error_u_vector10[109] + error_u_vector10[110] + error_u_vector10[111] + error_u_vector10[112] + error_u_vector10[113] + error_u_vector10[114] + error_u_vector10[115] + error_u_vector10[116] + error_u_vector10[117] + error_u_vector10[118] + error_u_vector10[119] + error_u_vector10[120] + error_u_vector10[121] + error_u_vector10[122] + error_u_vector10[123] + error_u_vector10[124] + error_u_vector10[125] + error_u_vector10[126] + error_u_vector10[127] + error_u_vector10[128] + error_u_vector10[129] + error_u_vector10[130] + error_u_vector10[131] + error_u_vector10[132] + error_u_vector10[133] + error_u_vector10[134] + error_u_vector10[135] + error_u_vector10[136] + error_u_vector10[137] + error_u_vector10[138] + error_u_vector10[139] + error_u_vector10[140] + error_u_vector10[141] + error_u_vector10[142] + error_u_vector10[143] + error_u_vector10[144] + error_u_vector10[145] + error_u_vector10[146] + error_u_vector10[147] + error_u_vector10[148] + error_u_vector10[149] + error_u_vector10[150] + error_u_vector10[151] + error_u_vector10[152] + error_u_vector10[153] + error_u_vector10[154] + error_u_vector10[155] + error_u_vector10[156] + error_u_vector10[157] + error_u_vector10[158] + error_u_vector10[159] + error_u_vector10[160] + error_u_vector10[161] + error_u_vector10[162] + error_u_vector10[163] + error_u_vector10[164] + error_u_vector10[165] + error_u_vector10[166] + error_u_vector10[167] + error_u_vector10[168] + error_u_vector10[169] + error_u_vector10[170] + error_u_vector10[171] + error_u_vector10[172] + error_u_vector10[173] + error_u_vector10[174] + error_u_vector10[175] + error_u_vector10[176] + error_u_vector10[177] + error_u_vector10[178] + error_u_vector10[179] + error_u_vector10[180] + error_u_vector10[181] + error_u_vector10[182] + error_u_vector10[183] + error_u_vector10[184] + error_u_vector10[185] + error_u_vector10[186] + error_u_vector10[187] + error_u_vector10[188] + error_u_vector10[189] + error_u_vector10[190] + error_u_vector10[191] + error_u_vector10[192] + error_u_vector10[193] + error_u_vector10[194] + error_u_vector10[195] + error_u_vector10[196] + error_u_vector10[197] + error_u_vector10[198] + error_u_vector10[199] + error_u_vector10[200] + error_u_vector10[201] + error_u_vector10[202] + error_u_vector10[203] + error_u_vector10[204] + error_u_vector10[205] + error_u_vector10[206] + error_u_vector10[207] + error_u_vector10[208] + error_u_vector10[209] + error_u_vector10[210] + error_u_vector10[211] + error_u_vector10[212] + error_u_vector10[213] + error_u_vector10[214] + error_u_vector10[215] + error_u_vector10[216] + error_u_vector10[217] + error_u_vector10[218] + error_u_vector10[219] + error_u_vector10[220] + error_u_vector10[221] + error_u_vector10[222] + error_u_vector10[223] + error_u_vector10[224] + error_u_vector10[225] + error_u_vector10[226] + error_u_vector10[227] + error_u_vector10[228] + error_u_vector10[229] + error_u_vector10[230] + error_u_vector10[231] + error_u_vector10[232] + error_u_vector10[233] + error_u_vector10[234] + error_u_vector10[235] + error_u_vector10[236] + error_u_vector10[237] + error_u_vector10[238]; 
            errs11_u <= error_u_vector11[0] + error_u_vector11[1] + error_u_vector11[2] + error_u_vector11[3] + error_u_vector11[4] + error_u_vector11[5] + error_u_vector11[6] + error_u_vector11[7] + error_u_vector11[8] + error_u_vector11[9] + error_u_vector11[10] + error_u_vector11[11] + error_u_vector11[12] + error_u_vector11[13] + error_u_vector11[14] + error_u_vector11[15] + error_u_vector11[16] + error_u_vector11[17] + error_u_vector11[18] + error_u_vector11[19] + error_u_vector11[20] + error_u_vector11[21] + error_u_vector11[22] + error_u_vector11[23] + error_u_vector11[24] + error_u_vector11[25] + error_u_vector11[26] + error_u_vector11[27] + error_u_vector11[28] + error_u_vector11[29] + error_u_vector11[30] + error_u_vector11[31] + error_u_vector11[32] + error_u_vector11[33] + error_u_vector11[34] + error_u_vector11[35] + error_u_vector11[36] + error_u_vector11[37] + error_u_vector11[38] + error_u_vector11[39] + error_u_vector11[40] + error_u_vector11[41] + error_u_vector11[42] + error_u_vector11[43] + error_u_vector11[44] + error_u_vector11[45] + error_u_vector11[46] + error_u_vector11[47] + error_u_vector11[48] + error_u_vector11[49] + error_u_vector11[50] + error_u_vector11[51] + error_u_vector11[52] + error_u_vector11[53] + error_u_vector11[54] + error_u_vector11[55] + error_u_vector11[56] + error_u_vector11[57] + error_u_vector11[58] + error_u_vector11[59] + error_u_vector11[60] + error_u_vector11[61] + error_u_vector11[62] + error_u_vector11[63] + error_u_vector11[64] + error_u_vector11[65] + error_u_vector11[66] + error_u_vector11[67] + error_u_vector11[68] + error_u_vector11[69] + error_u_vector11[70] + error_u_vector11[71] + error_u_vector11[72] + error_u_vector11[73] + error_u_vector11[74] + error_u_vector11[75] + error_u_vector11[76] + error_u_vector11[77] + error_u_vector11[78] + error_u_vector11[79] + error_u_vector11[80] + error_u_vector11[81] + error_u_vector11[82] + error_u_vector11[83] + error_u_vector11[84] + error_u_vector11[85] + error_u_vector11[86] + error_u_vector11[87] + error_u_vector11[88] + error_u_vector11[89] + error_u_vector11[90] + error_u_vector11[91] + error_u_vector11[92] + error_u_vector11[93] + error_u_vector11[94] + error_u_vector11[95] + error_u_vector11[96] + error_u_vector11[97] + error_u_vector11[98] + error_u_vector11[99] + error_u_vector11[100] + error_u_vector11[101] + error_u_vector11[102] + error_u_vector11[103] + error_u_vector11[104] + error_u_vector11[105] + error_u_vector11[106] + error_u_vector11[107] + error_u_vector11[108] + error_u_vector11[109] + error_u_vector11[110] + error_u_vector11[111] + error_u_vector11[112] + error_u_vector11[113] + error_u_vector11[114] + error_u_vector11[115] + error_u_vector11[116] + error_u_vector11[117] + error_u_vector11[118] + error_u_vector11[119] + error_u_vector11[120] + error_u_vector11[121] + error_u_vector11[122] + error_u_vector11[123] + error_u_vector11[124] + error_u_vector11[125] + error_u_vector11[126] + error_u_vector11[127] + error_u_vector11[128] + error_u_vector11[129] + error_u_vector11[130] + error_u_vector11[131] + error_u_vector11[132] + error_u_vector11[133] + error_u_vector11[134] + error_u_vector11[135] + error_u_vector11[136] + error_u_vector11[137] + error_u_vector11[138] + error_u_vector11[139] + error_u_vector11[140] + error_u_vector11[141] + error_u_vector11[142] + error_u_vector11[143] + error_u_vector11[144] + error_u_vector11[145] + error_u_vector11[146] + error_u_vector11[147] + error_u_vector11[148] + error_u_vector11[149] + error_u_vector11[150] + error_u_vector11[151] + error_u_vector11[152] + error_u_vector11[153] + error_u_vector11[154] + error_u_vector11[155] + error_u_vector11[156] + error_u_vector11[157] + error_u_vector11[158] + error_u_vector11[159] + error_u_vector11[160] + error_u_vector11[161] + error_u_vector11[162] + error_u_vector11[163] + error_u_vector11[164] + error_u_vector11[165] + error_u_vector11[166] + error_u_vector11[167] + error_u_vector11[168] + error_u_vector11[169] + error_u_vector11[170] + error_u_vector11[171] + error_u_vector11[172] + error_u_vector11[173] + error_u_vector11[174] + error_u_vector11[175] + error_u_vector11[176] + error_u_vector11[177] + error_u_vector11[178] + error_u_vector11[179] + error_u_vector11[180] + error_u_vector11[181] + error_u_vector11[182] + error_u_vector11[183] + error_u_vector11[184] + error_u_vector11[185] + error_u_vector11[186] + error_u_vector11[187] + error_u_vector11[188] + error_u_vector11[189] + error_u_vector11[190] + error_u_vector11[191] + error_u_vector11[192] + error_u_vector11[193] + error_u_vector11[194] + error_u_vector11[195] + error_u_vector11[196] + error_u_vector11[197] + error_u_vector11[198] + error_u_vector11[199] + error_u_vector11[200] + error_u_vector11[201] + error_u_vector11[202] + error_u_vector11[203] + error_u_vector11[204] + error_u_vector11[205] + error_u_vector11[206] + error_u_vector11[207] + error_u_vector11[208] + error_u_vector11[209] + error_u_vector11[210] + error_u_vector11[211] + error_u_vector11[212] + error_u_vector11[213] + error_u_vector11[214] + error_u_vector11[215] + error_u_vector11[216] + error_u_vector11[217] + error_u_vector11[218] + error_u_vector11[219] + error_u_vector11[220] + error_u_vector11[221] + error_u_vector11[222] + error_u_vector11[223] + error_u_vector11[224] + error_u_vector11[225] + error_u_vector11[226] + error_u_vector11[227] + error_u_vector11[228] + error_u_vector11[229] + error_u_vector11[230] + error_u_vector11[231] + error_u_vector11[232] + error_u_vector11[233] + error_u_vector11[234] + error_u_vector11[235] + error_u_vector11[236] + error_u_vector11[237] + error_u_vector11[238]; 
            errs12_u <= error_u_vector12[0] + error_u_vector12[1] + error_u_vector12[2] + error_u_vector12[3] + error_u_vector12[4] + error_u_vector12[5] + error_u_vector12[6] + error_u_vector12[7] + error_u_vector12[8] + error_u_vector12[9] + error_u_vector12[10] + error_u_vector12[11] + error_u_vector12[12] + error_u_vector12[13] + error_u_vector12[14] + error_u_vector12[15] + error_u_vector12[16] + error_u_vector12[17] + error_u_vector12[18] + error_u_vector12[19] + error_u_vector12[20] + error_u_vector12[21] + error_u_vector12[22] + error_u_vector12[23] + error_u_vector12[24] + error_u_vector12[25] + error_u_vector12[26] + error_u_vector12[27] + error_u_vector12[28] + error_u_vector12[29] + error_u_vector12[30] + error_u_vector12[31] + error_u_vector12[32] + error_u_vector12[33] + error_u_vector12[34] + error_u_vector12[35] + error_u_vector12[36] + error_u_vector12[37] + error_u_vector12[38] + error_u_vector12[39] + error_u_vector12[40] + error_u_vector12[41] + error_u_vector12[42] + error_u_vector12[43] + error_u_vector12[44] + error_u_vector12[45] + error_u_vector12[46] + error_u_vector12[47] + error_u_vector12[48] + error_u_vector12[49] + error_u_vector12[50] + error_u_vector12[51] + error_u_vector12[52] + error_u_vector12[53] + error_u_vector12[54] + error_u_vector12[55] + error_u_vector12[56] + error_u_vector12[57] + error_u_vector12[58] + error_u_vector12[59] + error_u_vector12[60] + error_u_vector12[61] + error_u_vector12[62] + error_u_vector12[63] + error_u_vector12[64] + error_u_vector12[65] + error_u_vector12[66] + error_u_vector12[67] + error_u_vector12[68] + error_u_vector12[69] + error_u_vector12[70] + error_u_vector12[71] + error_u_vector12[72] + error_u_vector12[73] + error_u_vector12[74] + error_u_vector12[75] + error_u_vector12[76] + error_u_vector12[77] + error_u_vector12[78] + error_u_vector12[79] + error_u_vector12[80] + error_u_vector12[81] + error_u_vector12[82] + error_u_vector12[83] + error_u_vector12[84] + error_u_vector12[85] + error_u_vector12[86] + error_u_vector12[87] + error_u_vector12[88] + error_u_vector12[89] + error_u_vector12[90] + error_u_vector12[91] + error_u_vector12[92] + error_u_vector12[93] + error_u_vector12[94] + error_u_vector12[95] + error_u_vector12[96] + error_u_vector12[97] + error_u_vector12[98] + error_u_vector12[99] + error_u_vector12[100] + error_u_vector12[101] + error_u_vector12[102] + error_u_vector12[103] + error_u_vector12[104] + error_u_vector12[105] + error_u_vector12[106] + error_u_vector12[107] + error_u_vector12[108] + error_u_vector12[109] + error_u_vector12[110] + error_u_vector12[111] + error_u_vector12[112] + error_u_vector12[113] + error_u_vector12[114] + error_u_vector12[115] + error_u_vector12[116] + error_u_vector12[117] + error_u_vector12[118] + error_u_vector12[119] + error_u_vector12[120] + error_u_vector12[121] + error_u_vector12[122] + error_u_vector12[123] + error_u_vector12[124] + error_u_vector12[125] + error_u_vector12[126] + error_u_vector12[127] + error_u_vector12[128] + error_u_vector12[129] + error_u_vector12[130] + error_u_vector12[131] + error_u_vector12[132] + error_u_vector12[133] + error_u_vector12[134] + error_u_vector12[135] + error_u_vector12[136] + error_u_vector12[137] + error_u_vector12[138] + error_u_vector12[139] + error_u_vector12[140] + error_u_vector12[141] + error_u_vector12[142] + error_u_vector12[143] + error_u_vector12[144] + error_u_vector12[145] + error_u_vector12[146] + error_u_vector12[147] + error_u_vector12[148] + error_u_vector12[149] + error_u_vector12[150] + error_u_vector12[151] + error_u_vector12[152] + error_u_vector12[153] + error_u_vector12[154] + error_u_vector12[155] + error_u_vector12[156] + error_u_vector12[157] + error_u_vector12[158] + error_u_vector12[159] + error_u_vector12[160] + error_u_vector12[161] + error_u_vector12[162] + error_u_vector12[163] + error_u_vector12[164] + error_u_vector12[165] + error_u_vector12[166] + error_u_vector12[167] + error_u_vector12[168] + error_u_vector12[169] + error_u_vector12[170] + error_u_vector12[171] + error_u_vector12[172] + error_u_vector12[173] + error_u_vector12[174] + error_u_vector12[175] + error_u_vector12[176] + error_u_vector12[177] + error_u_vector12[178] + error_u_vector12[179] + error_u_vector12[180] + error_u_vector12[181] + error_u_vector12[182] + error_u_vector12[183] + error_u_vector12[184] + error_u_vector12[185] + error_u_vector12[186] + error_u_vector12[187] + error_u_vector12[188] + error_u_vector12[189] + error_u_vector12[190] + error_u_vector12[191] + error_u_vector12[192] + error_u_vector12[193] + error_u_vector12[194] + error_u_vector12[195] + error_u_vector12[196] + error_u_vector12[197] + error_u_vector12[198] + error_u_vector12[199] + error_u_vector12[200] + error_u_vector12[201] + error_u_vector12[202] + error_u_vector12[203] + error_u_vector12[204] + error_u_vector12[205] + error_u_vector12[206] + error_u_vector12[207] + error_u_vector12[208] + error_u_vector12[209] + error_u_vector12[210] + error_u_vector12[211] + error_u_vector12[212] + error_u_vector12[213] + error_u_vector12[214] + error_u_vector12[215] + error_u_vector12[216] + error_u_vector12[217] + error_u_vector12[218] + error_u_vector12[219] + error_u_vector12[220] + error_u_vector12[221] + error_u_vector12[222] + error_u_vector12[223] + error_u_vector12[224] + error_u_vector12[225] + error_u_vector12[226] + error_u_vector12[227] + error_u_vector12[228] + error_u_vector12[229] + error_u_vector12[230] + error_u_vector12[231] + error_u_vector12[232] + error_u_vector12[233] + error_u_vector12[234] + error_u_vector12[235] + error_u_vector12[236] + error_u_vector12[237] + error_u_vector12[238]; 
            errs13_u <= error_u_vector13[0] + error_u_vector13[1] + error_u_vector13[2] + error_u_vector13[3] + error_u_vector13[4] + error_u_vector13[5] + error_u_vector13[6] + error_u_vector13[7] + error_u_vector13[8] + error_u_vector13[9] + error_u_vector13[10] + error_u_vector13[11] + error_u_vector13[12] + error_u_vector13[13] + error_u_vector13[14] + error_u_vector13[15] + error_u_vector13[16] + error_u_vector13[17] + error_u_vector13[18] + error_u_vector13[19] + error_u_vector13[20] + error_u_vector13[21] + error_u_vector13[22] + error_u_vector13[23] + error_u_vector13[24] + error_u_vector13[25] + error_u_vector13[26] + error_u_vector13[27] + error_u_vector13[28] + error_u_vector13[29] + error_u_vector13[30] + error_u_vector13[31] + error_u_vector13[32] + error_u_vector13[33] + error_u_vector13[34] + error_u_vector13[35] + error_u_vector13[36] + error_u_vector13[37] + error_u_vector13[38] + error_u_vector13[39] + error_u_vector13[40] + error_u_vector13[41] + error_u_vector13[42] + error_u_vector13[43] + error_u_vector13[44] + error_u_vector13[45] + error_u_vector13[46] + error_u_vector13[47] + error_u_vector13[48] + error_u_vector13[49] + error_u_vector13[50] + error_u_vector13[51] + error_u_vector13[52] + error_u_vector13[53] + error_u_vector13[54] + error_u_vector13[55] + error_u_vector13[56] + error_u_vector13[57] + error_u_vector13[58] + error_u_vector13[59] + error_u_vector13[60] + error_u_vector13[61] + error_u_vector13[62] + error_u_vector13[63] + error_u_vector13[64] + error_u_vector13[65] + error_u_vector13[66] + error_u_vector13[67] + error_u_vector13[68] + error_u_vector13[69] + error_u_vector13[70] + error_u_vector13[71] + error_u_vector13[72] + error_u_vector13[73] + error_u_vector13[74] + error_u_vector13[75] + error_u_vector13[76] + error_u_vector13[77] + error_u_vector13[78] + error_u_vector13[79] + error_u_vector13[80] + error_u_vector13[81] + error_u_vector13[82] + error_u_vector13[83] + error_u_vector13[84] + error_u_vector13[85] + error_u_vector13[86] + error_u_vector13[87] + error_u_vector13[88] + error_u_vector13[89] + error_u_vector13[90] + error_u_vector13[91] + error_u_vector13[92] + error_u_vector13[93] + error_u_vector13[94] + error_u_vector13[95] + error_u_vector13[96] + error_u_vector13[97] + error_u_vector13[98] + error_u_vector13[99] + error_u_vector13[100] + error_u_vector13[101] + error_u_vector13[102] + error_u_vector13[103] + error_u_vector13[104] + error_u_vector13[105] + error_u_vector13[106] + error_u_vector13[107] + error_u_vector13[108] + error_u_vector13[109] + error_u_vector13[110] + error_u_vector13[111] + error_u_vector13[112] + error_u_vector13[113] + error_u_vector13[114] + error_u_vector13[115] + error_u_vector13[116] + error_u_vector13[117] + error_u_vector13[118] + error_u_vector13[119] + error_u_vector13[120] + error_u_vector13[121] + error_u_vector13[122] + error_u_vector13[123] + error_u_vector13[124] + error_u_vector13[125] + error_u_vector13[126] + error_u_vector13[127] + error_u_vector13[128] + error_u_vector13[129] + error_u_vector13[130] + error_u_vector13[131] + error_u_vector13[132] + error_u_vector13[133] + error_u_vector13[134] + error_u_vector13[135] + error_u_vector13[136] + error_u_vector13[137] + error_u_vector13[138] + error_u_vector13[139] + error_u_vector13[140] + error_u_vector13[141] + error_u_vector13[142] + error_u_vector13[143] + error_u_vector13[144] + error_u_vector13[145] + error_u_vector13[146] + error_u_vector13[147] + error_u_vector13[148] + error_u_vector13[149] + error_u_vector13[150] + error_u_vector13[151] + error_u_vector13[152] + error_u_vector13[153] + error_u_vector13[154] + error_u_vector13[155] + error_u_vector13[156] + error_u_vector13[157] + error_u_vector13[158] + error_u_vector13[159] + error_u_vector13[160] + error_u_vector13[161] + error_u_vector13[162] + error_u_vector13[163] + error_u_vector13[164] + error_u_vector13[165] + error_u_vector13[166] + error_u_vector13[167] + error_u_vector13[168] + error_u_vector13[169] + error_u_vector13[170] + error_u_vector13[171] + error_u_vector13[172] + error_u_vector13[173] + error_u_vector13[174] + error_u_vector13[175] + error_u_vector13[176] + error_u_vector13[177] + error_u_vector13[178] + error_u_vector13[179] + error_u_vector13[180] + error_u_vector13[181] + error_u_vector13[182] + error_u_vector13[183] + error_u_vector13[184] + error_u_vector13[185] + error_u_vector13[186] + error_u_vector13[187] + error_u_vector13[188] + error_u_vector13[189] + error_u_vector13[190] + error_u_vector13[191] + error_u_vector13[192] + error_u_vector13[193] + error_u_vector13[194] + error_u_vector13[195] + error_u_vector13[196] + error_u_vector13[197] + error_u_vector13[198] + error_u_vector13[199] + error_u_vector13[200] + error_u_vector13[201] + error_u_vector13[202] + error_u_vector13[203] + error_u_vector13[204] + error_u_vector13[205] + error_u_vector13[206] + error_u_vector13[207] + error_u_vector13[208] + error_u_vector13[209] + error_u_vector13[210] + error_u_vector13[211] + error_u_vector13[212] + error_u_vector13[213] + error_u_vector13[214] + error_u_vector13[215] + error_u_vector13[216] + error_u_vector13[217] + error_u_vector13[218] + error_u_vector13[219] + error_u_vector13[220] + error_u_vector13[221] + error_u_vector13[222] + error_u_vector13[223] + error_u_vector13[224] + error_u_vector13[225] + error_u_vector13[226] + error_u_vector13[227] + error_u_vector13[228] + error_u_vector13[229] + error_u_vector13[230] + error_u_vector13[231] + error_u_vector13[232] + error_u_vector13[233] + error_u_vector13[234] + error_u_vector13[235] + error_u_vector13[236] + error_u_vector13[237] + error_u_vector13[238]; 
            errs14_u <= error_u_vector14[0] + error_u_vector14[1] + error_u_vector14[2] + error_u_vector14[3] + error_u_vector14[4] + error_u_vector14[5] + error_u_vector14[6] + error_u_vector14[7] + error_u_vector14[8] + error_u_vector14[9] + error_u_vector14[10] + error_u_vector14[11] + error_u_vector14[12] + error_u_vector14[13] + error_u_vector14[14] + error_u_vector14[15] + error_u_vector14[16] + error_u_vector14[17] + error_u_vector14[18] + error_u_vector14[19] + error_u_vector14[20] + error_u_vector14[21] + error_u_vector14[22] + error_u_vector14[23] + error_u_vector14[24] + error_u_vector14[25] + error_u_vector14[26] + error_u_vector14[27] + error_u_vector14[28] + error_u_vector14[29] + error_u_vector14[30] + error_u_vector14[31] + error_u_vector14[32] + error_u_vector14[33] + error_u_vector14[34] + error_u_vector14[35] + error_u_vector14[36] + error_u_vector14[37] + error_u_vector14[38] + error_u_vector14[39] + error_u_vector14[40] + error_u_vector14[41] + error_u_vector14[42] + error_u_vector14[43] + error_u_vector14[44] + error_u_vector14[45] + error_u_vector14[46] + error_u_vector14[47] + error_u_vector14[48] + error_u_vector14[49] + error_u_vector14[50] + error_u_vector14[51] + error_u_vector14[52] + error_u_vector14[53] + error_u_vector14[54] + error_u_vector14[55] + error_u_vector14[56] + error_u_vector14[57] + error_u_vector14[58] + error_u_vector14[59] + error_u_vector14[60] + error_u_vector14[61] + error_u_vector14[62] + error_u_vector14[63] + error_u_vector14[64] + error_u_vector14[65] + error_u_vector14[66] + error_u_vector14[67] + error_u_vector14[68] + error_u_vector14[69] + error_u_vector14[70] + error_u_vector14[71] + error_u_vector14[72] + error_u_vector14[73] + error_u_vector14[74] + error_u_vector14[75] + error_u_vector14[76] + error_u_vector14[77] + error_u_vector14[78] + error_u_vector14[79] + error_u_vector14[80] + error_u_vector14[81] + error_u_vector14[82] + error_u_vector14[83] + error_u_vector14[84] + error_u_vector14[85] + error_u_vector14[86] + error_u_vector14[87] + error_u_vector14[88] + error_u_vector14[89] + error_u_vector14[90] + error_u_vector14[91] + error_u_vector14[92] + error_u_vector14[93] + error_u_vector14[94] + error_u_vector14[95] + error_u_vector14[96] + error_u_vector14[97] + error_u_vector14[98] + error_u_vector14[99] + error_u_vector14[100] + error_u_vector14[101] + error_u_vector14[102] + error_u_vector14[103] + error_u_vector14[104] + error_u_vector14[105] + error_u_vector14[106] + error_u_vector14[107] + error_u_vector14[108] + error_u_vector14[109] + error_u_vector14[110] + error_u_vector14[111] + error_u_vector14[112] + error_u_vector14[113] + error_u_vector14[114] + error_u_vector14[115] + error_u_vector14[116] + error_u_vector14[117] + error_u_vector14[118] + error_u_vector14[119] + error_u_vector14[120] + error_u_vector14[121] + error_u_vector14[122] + error_u_vector14[123] + error_u_vector14[124] + error_u_vector14[125] + error_u_vector14[126] + error_u_vector14[127] + error_u_vector14[128] + error_u_vector14[129] + error_u_vector14[130] + error_u_vector14[131] + error_u_vector14[132] + error_u_vector14[133] + error_u_vector14[134] + error_u_vector14[135] + error_u_vector14[136] + error_u_vector14[137] + error_u_vector14[138] + error_u_vector14[139] + error_u_vector14[140] + error_u_vector14[141] + error_u_vector14[142] + error_u_vector14[143] + error_u_vector14[144] + error_u_vector14[145] + error_u_vector14[146] + error_u_vector14[147] + error_u_vector14[148] + error_u_vector14[149] + error_u_vector14[150] + error_u_vector14[151] + error_u_vector14[152] + error_u_vector14[153] + error_u_vector14[154] + error_u_vector14[155] + error_u_vector14[156] + error_u_vector14[157] + error_u_vector14[158] + error_u_vector14[159] + error_u_vector14[160] + error_u_vector14[161] + error_u_vector14[162] + error_u_vector14[163] + error_u_vector14[164] + error_u_vector14[165] + error_u_vector14[166] + error_u_vector14[167] + error_u_vector14[168] + error_u_vector14[169] + error_u_vector14[170] + error_u_vector14[171] + error_u_vector14[172] + error_u_vector14[173] + error_u_vector14[174] + error_u_vector14[175] + error_u_vector14[176] + error_u_vector14[177] + error_u_vector14[178] + error_u_vector14[179] + error_u_vector14[180] + error_u_vector14[181] + error_u_vector14[182] + error_u_vector14[183] + error_u_vector14[184] + error_u_vector14[185] + error_u_vector14[186] + error_u_vector14[187] + error_u_vector14[188] + error_u_vector14[189] + error_u_vector14[190] + error_u_vector14[191] + error_u_vector14[192] + error_u_vector14[193] + error_u_vector14[194] + error_u_vector14[195] + error_u_vector14[196] + error_u_vector14[197] + error_u_vector14[198] + error_u_vector14[199] + error_u_vector14[200] + error_u_vector14[201] + error_u_vector14[202] + error_u_vector14[203] + error_u_vector14[204] + error_u_vector14[205] + error_u_vector14[206] + error_u_vector14[207] + error_u_vector14[208] + error_u_vector14[209] + error_u_vector14[210] + error_u_vector14[211] + error_u_vector14[212] + error_u_vector14[213] + error_u_vector14[214] + error_u_vector14[215] + error_u_vector14[216] + error_u_vector14[217] + error_u_vector14[218] + error_u_vector14[219] + error_u_vector14[220] + error_u_vector14[221] + error_u_vector14[222] + error_u_vector14[223] + error_u_vector14[224] + error_u_vector14[225] + error_u_vector14[226] + error_u_vector14[227] + error_u_vector14[228] + error_u_vector14[229] + error_u_vector14[230] + error_u_vector14[231] + error_u_vector14[232] + error_u_vector14[233] + error_u_vector14[234] + error_u_vector14[235] + error_u_vector14[236] + error_u_vector14[237] + error_u_vector14[238]; 
            errs15_u <= error_u_vector15[0] + error_u_vector15[1] + error_u_vector15[2] + error_u_vector15[3] + error_u_vector15[4] + error_u_vector15[5] + error_u_vector15[6] + error_u_vector15[7] + error_u_vector15[8] + error_u_vector15[9] + error_u_vector15[10] + error_u_vector15[11] + error_u_vector15[12] + error_u_vector15[13] + error_u_vector15[14] + error_u_vector15[15] + error_u_vector15[16] + error_u_vector15[17] + error_u_vector15[18] + error_u_vector15[19] + error_u_vector15[20] + error_u_vector15[21] + error_u_vector15[22] + error_u_vector15[23] + error_u_vector15[24] + error_u_vector15[25] + error_u_vector15[26] + error_u_vector15[27] + error_u_vector15[28] + error_u_vector15[29] + error_u_vector15[30] + error_u_vector15[31] + error_u_vector15[32] + error_u_vector15[33] + error_u_vector15[34] + error_u_vector15[35] + error_u_vector15[36] + error_u_vector15[37] + error_u_vector15[38] + error_u_vector15[39] + error_u_vector15[40] + error_u_vector15[41] + error_u_vector15[42] + error_u_vector15[43] + error_u_vector15[44] + error_u_vector15[45] + error_u_vector15[46] + error_u_vector15[47] + error_u_vector15[48] + error_u_vector15[49] + error_u_vector15[50] + error_u_vector15[51] + error_u_vector15[52] + error_u_vector15[53] + error_u_vector15[54] + error_u_vector15[55] + error_u_vector15[56] + error_u_vector15[57] + error_u_vector15[58] + error_u_vector15[59] + error_u_vector15[60] + error_u_vector15[61] + error_u_vector15[62] + error_u_vector15[63] + error_u_vector15[64] + error_u_vector15[65] + error_u_vector15[66] + error_u_vector15[67] + error_u_vector15[68] + error_u_vector15[69] + error_u_vector15[70] + error_u_vector15[71] + error_u_vector15[72] + error_u_vector15[73] + error_u_vector15[74] + error_u_vector15[75] + error_u_vector15[76] + error_u_vector15[77] + error_u_vector15[78] + error_u_vector15[79] + error_u_vector15[80] + error_u_vector15[81] + error_u_vector15[82] + error_u_vector15[83] + error_u_vector15[84] + error_u_vector15[85] + error_u_vector15[86] + error_u_vector15[87] + error_u_vector15[88] + error_u_vector15[89] + error_u_vector15[90] + error_u_vector15[91] + error_u_vector15[92] + error_u_vector15[93] + error_u_vector15[94] + error_u_vector15[95] + error_u_vector15[96] + error_u_vector15[97] + error_u_vector15[98] + error_u_vector15[99] + error_u_vector15[100] + error_u_vector15[101] + error_u_vector15[102] + error_u_vector15[103] + error_u_vector15[104] + error_u_vector15[105] + error_u_vector15[106] + error_u_vector15[107] + error_u_vector15[108] + error_u_vector15[109] + error_u_vector15[110] + error_u_vector15[111] + error_u_vector15[112] + error_u_vector15[113] + error_u_vector15[114] + error_u_vector15[115] + error_u_vector15[116] + error_u_vector15[117] + error_u_vector15[118] + error_u_vector15[119] + error_u_vector15[120] + error_u_vector15[121] + error_u_vector15[122] + error_u_vector15[123] + error_u_vector15[124] + error_u_vector15[125] + error_u_vector15[126] + error_u_vector15[127] + error_u_vector15[128] + error_u_vector15[129] + error_u_vector15[130] + error_u_vector15[131] + error_u_vector15[132] + error_u_vector15[133] + error_u_vector15[134] + error_u_vector15[135] + error_u_vector15[136] + error_u_vector15[137] + error_u_vector15[138] + error_u_vector15[139] + error_u_vector15[140] + error_u_vector15[141] + error_u_vector15[142] + error_u_vector15[143] + error_u_vector15[144] + error_u_vector15[145] + error_u_vector15[146] + error_u_vector15[147] + error_u_vector15[148] + error_u_vector15[149] + error_u_vector15[150] + error_u_vector15[151] + error_u_vector15[152] + error_u_vector15[153] + error_u_vector15[154] + error_u_vector15[155] + error_u_vector15[156] + error_u_vector15[157] + error_u_vector15[158] + error_u_vector15[159] + error_u_vector15[160] + error_u_vector15[161] + error_u_vector15[162] + error_u_vector15[163] + error_u_vector15[164] + error_u_vector15[165] + error_u_vector15[166] + error_u_vector15[167] + error_u_vector15[168] + error_u_vector15[169] + error_u_vector15[170] + error_u_vector15[171] + error_u_vector15[172] + error_u_vector15[173] + error_u_vector15[174] + error_u_vector15[175] + error_u_vector15[176] + error_u_vector15[177] + error_u_vector15[178] + error_u_vector15[179] + error_u_vector15[180] + error_u_vector15[181] + error_u_vector15[182] + error_u_vector15[183] + error_u_vector15[184] + error_u_vector15[185] + error_u_vector15[186] + error_u_vector15[187] + error_u_vector15[188] + error_u_vector15[189] + error_u_vector15[190] + error_u_vector15[191] + error_u_vector15[192] + error_u_vector15[193] + error_u_vector15[194] + error_u_vector15[195] + error_u_vector15[196] + error_u_vector15[197] + error_u_vector15[198] + error_u_vector15[199] + error_u_vector15[200] + error_u_vector15[201] + error_u_vector15[202] + error_u_vector15[203] + error_u_vector15[204] + error_u_vector15[205] + error_u_vector15[206] + error_u_vector15[207] + error_u_vector15[208] + error_u_vector15[209] + error_u_vector15[210] + error_u_vector15[211] + error_u_vector15[212] + error_u_vector15[213] + error_u_vector15[214] + error_u_vector15[215] + error_u_vector15[216] + error_u_vector15[217] + error_u_vector15[218] + error_u_vector15[219] + error_u_vector15[220] + error_u_vector15[221] + error_u_vector15[222] + error_u_vector15[223] + error_u_vector15[224] + error_u_vector15[225] + error_u_vector15[226] + error_u_vector15[227] + error_u_vector15[228] + error_u_vector15[229] + error_u_vector15[230] + error_u_vector15[231] + error_u_vector15[232] + error_u_vector15[233] + error_u_vector15[234] + error_u_vector15[235] + error_u_vector15[236] + error_u_vector15[237] + error_u_vector15[238]; 
            errs16_u <= error_u_vector16[0] + error_u_vector16[1] + error_u_vector16[2] + error_u_vector16[3] + error_u_vector16[4] + error_u_vector16[5] + error_u_vector16[6] + error_u_vector16[7] + error_u_vector16[8] + error_u_vector16[9] + error_u_vector16[10] + error_u_vector16[11] + error_u_vector16[12] + error_u_vector16[13] + error_u_vector16[14] + error_u_vector16[15] + error_u_vector16[16] + error_u_vector16[17] + error_u_vector16[18] + error_u_vector16[19] + error_u_vector16[20] + error_u_vector16[21] + error_u_vector16[22] + error_u_vector16[23] + error_u_vector16[24] + error_u_vector16[25] + error_u_vector16[26] + error_u_vector16[27] + error_u_vector16[28] + error_u_vector16[29] + error_u_vector16[30] + error_u_vector16[31] + error_u_vector16[32] + error_u_vector16[33] + error_u_vector16[34] + error_u_vector16[35] + error_u_vector16[36] + error_u_vector16[37] + error_u_vector16[38] + error_u_vector16[39] + error_u_vector16[40] + error_u_vector16[41] + error_u_vector16[42] + error_u_vector16[43] + error_u_vector16[44] + error_u_vector16[45] + error_u_vector16[46] + error_u_vector16[47] + error_u_vector16[48] + error_u_vector16[49] + error_u_vector16[50] + error_u_vector16[51] + error_u_vector16[52] + error_u_vector16[53] + error_u_vector16[54] + error_u_vector16[55] + error_u_vector16[56] + error_u_vector16[57] + error_u_vector16[58] + error_u_vector16[59] + error_u_vector16[60] + error_u_vector16[61] + error_u_vector16[62] + error_u_vector16[63] + error_u_vector16[64] + error_u_vector16[65] + error_u_vector16[66] + error_u_vector16[67] + error_u_vector16[68] + error_u_vector16[69] + error_u_vector16[70] + error_u_vector16[71] + error_u_vector16[72] + error_u_vector16[73] + error_u_vector16[74] + error_u_vector16[75] + error_u_vector16[76] + error_u_vector16[77] + error_u_vector16[78] + error_u_vector16[79] + error_u_vector16[80] + error_u_vector16[81] + error_u_vector16[82] + error_u_vector16[83] + error_u_vector16[84] + error_u_vector16[85] + error_u_vector16[86] + error_u_vector16[87] + error_u_vector16[88] + error_u_vector16[89] + error_u_vector16[90] + error_u_vector16[91] + error_u_vector16[92] + error_u_vector16[93] + error_u_vector16[94] + error_u_vector16[95] + error_u_vector16[96] + error_u_vector16[97] + error_u_vector16[98] + error_u_vector16[99] + error_u_vector16[100] + error_u_vector16[101] + error_u_vector16[102] + error_u_vector16[103] + error_u_vector16[104] + error_u_vector16[105] + error_u_vector16[106] + error_u_vector16[107] + error_u_vector16[108] + error_u_vector16[109] + error_u_vector16[110] + error_u_vector16[111] + error_u_vector16[112] + error_u_vector16[113] + error_u_vector16[114] + error_u_vector16[115] + error_u_vector16[116] + error_u_vector16[117] + error_u_vector16[118] + error_u_vector16[119] + error_u_vector16[120] + error_u_vector16[121] + error_u_vector16[122] + error_u_vector16[123] + error_u_vector16[124] + error_u_vector16[125] + error_u_vector16[126] + error_u_vector16[127] + error_u_vector16[128] + error_u_vector16[129] + error_u_vector16[130] + error_u_vector16[131] + error_u_vector16[132] + error_u_vector16[133] + error_u_vector16[134] + error_u_vector16[135] + error_u_vector16[136] + error_u_vector16[137] + error_u_vector16[138] + error_u_vector16[139] + error_u_vector16[140] + error_u_vector16[141] + error_u_vector16[142] + error_u_vector16[143] + error_u_vector16[144] + error_u_vector16[145] + error_u_vector16[146] + error_u_vector16[147] + error_u_vector16[148] + error_u_vector16[149] + error_u_vector16[150] + error_u_vector16[151] + error_u_vector16[152] + error_u_vector16[153] + error_u_vector16[154] + error_u_vector16[155] + error_u_vector16[156] + error_u_vector16[157] + error_u_vector16[158] + error_u_vector16[159] + error_u_vector16[160] + error_u_vector16[161] + error_u_vector16[162] + error_u_vector16[163] + error_u_vector16[164] + error_u_vector16[165] + error_u_vector16[166] + error_u_vector16[167] + error_u_vector16[168] + error_u_vector16[169] + error_u_vector16[170] + error_u_vector16[171] + error_u_vector16[172] + error_u_vector16[173] + error_u_vector16[174] + error_u_vector16[175] + error_u_vector16[176] + error_u_vector16[177] + error_u_vector16[178] + error_u_vector16[179] + error_u_vector16[180] + error_u_vector16[181] + error_u_vector16[182] + error_u_vector16[183] + error_u_vector16[184] + error_u_vector16[185] + error_u_vector16[186] + error_u_vector16[187] + error_u_vector16[188] + error_u_vector16[189] + error_u_vector16[190] + error_u_vector16[191] + error_u_vector16[192] + error_u_vector16[193] + error_u_vector16[194] + error_u_vector16[195] + error_u_vector16[196] + error_u_vector16[197] + error_u_vector16[198] + error_u_vector16[199] + error_u_vector16[200] + error_u_vector16[201] + error_u_vector16[202] + error_u_vector16[203] + error_u_vector16[204] + error_u_vector16[205] + error_u_vector16[206] + error_u_vector16[207] + error_u_vector16[208] + error_u_vector16[209] + error_u_vector16[210] + error_u_vector16[211] + error_u_vector16[212] + error_u_vector16[213] + error_u_vector16[214] + error_u_vector16[215] + error_u_vector16[216] + error_u_vector16[217] + error_u_vector16[218] + error_u_vector16[219] + error_u_vector16[220] + error_u_vector16[221] + error_u_vector16[222] + error_u_vector16[223] + error_u_vector16[224] + error_u_vector16[225] + error_u_vector16[226] + error_u_vector16[227] + error_u_vector16[228] + error_u_vector16[229] + error_u_vector16[230] + error_u_vector16[231] + error_u_vector16[232] + error_u_vector16[233] + error_u_vector16[234] + error_u_vector16[235] + error_u_vector16[236] + error_u_vector16[237] + error_u_vector16[238]; 
  
            errs1 <= error_vector1[0] + error_vector1[1] + error_vector1[2] + error_vector1[3] + error_vector1[4] + error_vector1[5] + error_vector1[6] + error_vector1[7] + error_vector1[8] + error_vector1[9] + error_vector1[10] + error_vector1[11] + error_vector1[12] + error_vector1[13] + error_vector1[14] + error_vector1[15] + error_vector1[16] + error_vector1[17] + error_vector1[18] + error_vector1[19] + error_vector1[20] + error_vector1[21] + error_vector1[22] + error_vector1[23] + error_vector1[24] + error_vector1[25] + error_vector1[26] + error_vector1[27] + error_vector1[28] + error_vector1[29] + error_vector1[30] + error_vector1[31] + error_vector1[32] + error_vector1[33] + error_vector1[34] + error_vector1[35] + error_vector1[36] + error_vector1[37] + error_vector1[38] + error_vector1[39] + error_vector1[40] + error_vector1[41] + error_vector1[42] + error_vector1[43] + error_vector1[44] + error_vector1[45] + error_vector1[46] + error_vector1[47] + error_vector1[48] + error_vector1[49] + error_vector1[50] + error_vector1[51] + error_vector1[52] + error_vector1[53] + error_vector1[54] + error_vector1[55] + error_vector1[56] + error_vector1[57] + error_vector1[58] + error_vector1[59] + error_vector1[60] + error_vector1[61] + error_vector1[62] + error_vector1[63] + error_vector1[64] + error_vector1[65] + error_vector1[66] + error_vector1[67] + error_vector1[68] + error_vector1[69] + error_vector1[70] + error_vector1[71] + error_vector1[72] + error_vector1[73] + error_vector1[74] + error_vector1[75] + error_vector1[76] + error_vector1[77] + error_vector1[78] + error_vector1[79] + error_vector1[80] + error_vector1[81] + error_vector1[82] + error_vector1[83] + error_vector1[84] + error_vector1[85] + error_vector1[86] + error_vector1[87] + error_vector1[88] + error_vector1[89] + error_vector1[90] + error_vector1[91] + error_vector1[92] + error_vector1[93] + error_vector1[94] + error_vector1[95] + error_vector1[96] + error_vector1[97] + error_vector1[98] + error_vector1[99] + error_vector1[100] + error_vector1[101] + error_vector1[102] + error_vector1[103] + error_vector1[104] + error_vector1[105] + error_vector1[106] + error_vector1[107] + error_vector1[108] + error_vector1[109] + error_vector1[110] + error_vector1[111] + error_vector1[112] + error_vector1[113] + error_vector1[114] + error_vector1[115] + error_vector1[116] + error_vector1[117] + error_vector1[118] + error_vector1[119] + error_vector1[120] + error_vector1[121] + error_vector1[122] + error_vector1[123] + error_vector1[124] + error_vector1[125] + error_vector1[126] + error_vector1[127] + error_vector1[128] + error_vector1[129] + error_vector1[130] + error_vector1[131] + error_vector1[132] + error_vector1[133] + error_vector1[134] + error_vector1[135] + error_vector1[136] + error_vector1[137] + error_vector1[138] + error_vector1[139] + error_vector1[140] + error_vector1[141] + error_vector1[142] + error_vector1[143] + error_vector1[144] + error_vector1[145] + error_vector1[146] + error_vector1[147] + error_vector1[148] + error_vector1[149] + error_vector1[150] + error_vector1[151] + error_vector1[152] + error_vector1[153] + error_vector1[154] + error_vector1[155] + error_vector1[156] + error_vector1[157] + error_vector1[158] + error_vector1[159] + error_vector1[160] + error_vector1[161] + error_vector1[162] + error_vector1[163] + error_vector1[164] + error_vector1[165] + error_vector1[166] + error_vector1[167] + error_vector1[168] + error_vector1[169] + error_vector1[170] + error_vector1[171] + error_vector1[172] + error_vector1[173] + error_vector1[174] + error_vector1[175] + error_vector1[176] + error_vector1[177] + error_vector1[178] + error_vector1[179] + error_vector1[180] + error_vector1[181] + error_vector1[182] + error_vector1[183] + error_vector1[184] + error_vector1[185] + error_vector1[186] + error_vector1[187] + error_vector1[188] + error_vector1[189] + error_vector1[190] + error_vector1[191] + error_vector1[192] + error_vector1[193] + error_vector1[194] + error_vector1[195] + error_vector1[196] + error_vector1[197] + error_vector1[198] + error_vector1[199] + error_vector1[200] + error_vector1[201] + error_vector1[202] + error_vector1[203] + error_vector1[204] + error_vector1[205] + error_vector1[206] + error_vector1[207] + error_vector1[208] + error_vector1[209] + error_vector1[210] + error_vector1[211] + error_vector1[212] + error_vector1[213] + error_vector1[214] + error_vector1[215] + error_vector1[216] + error_vector1[217] + error_vector1[218] + error_vector1[219] + error_vector1[220] + error_vector1[221] + error_vector1[222] + error_vector1[223] + error_vector1[224] + error_vector1[225] + error_vector1[226] + error_vector1[227] + error_vector1[228] + error_vector1[229] + error_vector1[230] + error_vector1[231] + error_vector1[232] + error_vector1[233] + error_vector1[234] + error_vector1[235] + error_vector1[236] + error_vector1[237] + error_vector1[238]; 
            errs2 <= error_vector2[0] + error_vector2[1] + error_vector2[2] + error_vector2[3] + error_vector2[4] + error_vector2[5] + error_vector2[6] + error_vector2[7] + error_vector2[8] + error_vector2[9] + error_vector2[10] + error_vector2[11] + error_vector2[12] + error_vector2[13] + error_vector2[14] + error_vector2[15] + error_vector2[16] + error_vector2[17] + error_vector2[18] + error_vector2[19] + error_vector2[20] + error_vector2[21] + error_vector2[22] + error_vector2[23] + error_vector2[24] + error_vector2[25] + error_vector2[26] + error_vector2[27] + error_vector2[28] + error_vector2[29] + error_vector2[30] + error_vector2[31] + error_vector2[32] + error_vector2[33] + error_vector2[34] + error_vector2[35] + error_vector2[36] + error_vector2[37] + error_vector2[38] + error_vector2[39] + error_vector2[40] + error_vector2[41] + error_vector2[42] + error_vector2[43] + error_vector2[44] + error_vector2[45] + error_vector2[46] + error_vector2[47] + error_vector2[48] + error_vector2[49] + error_vector2[50] + error_vector2[51] + error_vector2[52] + error_vector2[53] + error_vector2[54] + error_vector2[55] + error_vector2[56] + error_vector2[57] + error_vector2[58] + error_vector2[59] + error_vector2[60] + error_vector2[61] + error_vector2[62] + error_vector2[63] + error_vector2[64] + error_vector2[65] + error_vector2[66] + error_vector2[67] + error_vector2[68] + error_vector2[69] + error_vector2[70] + error_vector2[71] + error_vector2[72] + error_vector2[73] + error_vector2[74] + error_vector2[75] + error_vector2[76] + error_vector2[77] + error_vector2[78] + error_vector2[79] + error_vector2[80] + error_vector2[81] + error_vector2[82] + error_vector2[83] + error_vector2[84] + error_vector2[85] + error_vector2[86] + error_vector2[87] + error_vector2[88] + error_vector2[89] + error_vector2[90] + error_vector2[91] + error_vector2[92] + error_vector2[93] + error_vector2[94] + error_vector2[95] + error_vector2[96] + error_vector2[97] + error_vector2[98] + error_vector2[99] + error_vector2[100] + error_vector2[101] + error_vector2[102] + error_vector2[103] + error_vector2[104] + error_vector2[105] + error_vector2[106] + error_vector2[107] + error_vector2[108] + error_vector2[109] + error_vector2[110] + error_vector2[111] + error_vector2[112] + error_vector2[113] + error_vector2[114] + error_vector2[115] + error_vector2[116] + error_vector2[117] + error_vector2[118] + error_vector2[119] + error_vector2[120] + error_vector2[121] + error_vector2[122] + error_vector2[123] + error_vector2[124] + error_vector2[125] + error_vector2[126] + error_vector2[127] + error_vector2[128] + error_vector2[129] + error_vector2[130] + error_vector2[131] + error_vector2[132] + error_vector2[133] + error_vector2[134] + error_vector2[135] + error_vector2[136] + error_vector2[137] + error_vector2[138] + error_vector2[139] + error_vector2[140] + error_vector2[141] + error_vector2[142] + error_vector2[143] + error_vector2[144] + error_vector2[145] + error_vector2[146] + error_vector2[147] + error_vector2[148] + error_vector2[149] + error_vector2[150] + error_vector2[151] + error_vector2[152] + error_vector2[153] + error_vector2[154] + error_vector2[155] + error_vector2[156] + error_vector2[157] + error_vector2[158] + error_vector2[159] + error_vector2[160] + error_vector2[161] + error_vector2[162] + error_vector2[163] + error_vector2[164] + error_vector2[165] + error_vector2[166] + error_vector2[167] + error_vector2[168] + error_vector2[169] + error_vector2[170] + error_vector2[171] + error_vector2[172] + error_vector2[173] + error_vector2[174] + error_vector2[175] + error_vector2[176] + error_vector2[177] + error_vector2[178] + error_vector2[179] + error_vector2[180] + error_vector2[181] + error_vector2[182] + error_vector2[183] + error_vector2[184] + error_vector2[185] + error_vector2[186] + error_vector2[187] + error_vector2[188] + error_vector2[189] + error_vector2[190] + error_vector2[191] + error_vector2[192] + error_vector2[193] + error_vector2[194] + error_vector2[195] + error_vector2[196] + error_vector2[197] + error_vector2[198] + error_vector2[199] + error_vector2[200] + error_vector2[201] + error_vector2[202] + error_vector2[203] + error_vector2[204] + error_vector2[205] + error_vector2[206] + error_vector2[207] + error_vector2[208] + error_vector2[209] + error_vector2[210] + error_vector2[211] + error_vector2[212] + error_vector2[213] + error_vector2[214] + error_vector2[215] + error_vector2[216] + error_vector2[217] + error_vector2[218] + error_vector2[219] + error_vector2[220] + error_vector2[221] + error_vector2[222] + error_vector2[223] + error_vector2[224] + error_vector2[225] + error_vector2[226] + error_vector2[227] + error_vector2[228] + error_vector2[229] + error_vector2[230] + error_vector2[231] + error_vector2[232] + error_vector2[233] + error_vector2[234] + error_vector2[235] + error_vector2[236] + error_vector2[237] + error_vector2[238]; 
            errs3 <= error_vector3[0] + error_vector3[1] + error_vector3[2] + error_vector3[3] + error_vector3[4] + error_vector3[5] + error_vector3[6] + error_vector3[7] + error_vector3[8] + error_vector3[9] + error_vector3[10] + error_vector3[11] + error_vector3[12] + error_vector3[13] + error_vector3[14] + error_vector3[15] + error_vector3[16] + error_vector3[17] + error_vector3[18] + error_vector3[19] + error_vector3[20] + error_vector3[21] + error_vector3[22] + error_vector3[23] + error_vector3[24] + error_vector3[25] + error_vector3[26] + error_vector3[27] + error_vector3[28] + error_vector3[29] + error_vector3[30] + error_vector3[31] + error_vector3[32] + error_vector3[33] + error_vector3[34] + error_vector3[35] + error_vector3[36] + error_vector3[37] + error_vector3[38] + error_vector3[39] + error_vector3[40] + error_vector3[41] + error_vector3[42] + error_vector3[43] + error_vector3[44] + error_vector3[45] + error_vector3[46] + error_vector3[47] + error_vector3[48] + error_vector3[49] + error_vector3[50] + error_vector3[51] + error_vector3[52] + error_vector3[53] + error_vector3[54] + error_vector3[55] + error_vector3[56] + error_vector3[57] + error_vector3[58] + error_vector3[59] + error_vector3[60] + error_vector3[61] + error_vector3[62] + error_vector3[63] + error_vector3[64] + error_vector3[65] + error_vector3[66] + error_vector3[67] + error_vector3[68] + error_vector3[69] + error_vector3[70] + error_vector3[71] + error_vector3[72] + error_vector3[73] + error_vector3[74] + error_vector3[75] + error_vector3[76] + error_vector3[77] + error_vector3[78] + error_vector3[79] + error_vector3[80] + error_vector3[81] + error_vector3[82] + error_vector3[83] + error_vector3[84] + error_vector3[85] + error_vector3[86] + error_vector3[87] + error_vector3[88] + error_vector3[89] + error_vector3[90] + error_vector3[91] + error_vector3[92] + error_vector3[93] + error_vector3[94] + error_vector3[95] + error_vector3[96] + error_vector3[97] + error_vector3[98] + error_vector3[99] + error_vector3[100] + error_vector3[101] + error_vector3[102] + error_vector3[103] + error_vector3[104] + error_vector3[105] + error_vector3[106] + error_vector3[107] + error_vector3[108] + error_vector3[109] + error_vector3[110] + error_vector3[111] + error_vector3[112] + error_vector3[113] + error_vector3[114] + error_vector3[115] + error_vector3[116] + error_vector3[117] + error_vector3[118] + error_vector3[119] + error_vector3[120] + error_vector3[121] + error_vector3[122] + error_vector3[123] + error_vector3[124] + error_vector3[125] + error_vector3[126] + error_vector3[127] + error_vector3[128] + error_vector3[129] + error_vector3[130] + error_vector3[131] + error_vector3[132] + error_vector3[133] + error_vector3[134] + error_vector3[135] + error_vector3[136] + error_vector3[137] + error_vector3[138] + error_vector3[139] + error_vector3[140] + error_vector3[141] + error_vector3[142] + error_vector3[143] + error_vector3[144] + error_vector3[145] + error_vector3[146] + error_vector3[147] + error_vector3[148] + error_vector3[149] + error_vector3[150] + error_vector3[151] + error_vector3[152] + error_vector3[153] + error_vector3[154] + error_vector3[155] + error_vector3[156] + error_vector3[157] + error_vector3[158] + error_vector3[159] + error_vector3[160] + error_vector3[161] + error_vector3[162] + error_vector3[163] + error_vector3[164] + error_vector3[165] + error_vector3[166] + error_vector3[167] + error_vector3[168] + error_vector3[169] + error_vector3[170] + error_vector3[171] + error_vector3[172] + error_vector3[173] + error_vector3[174] + error_vector3[175] + error_vector3[176] + error_vector3[177] + error_vector3[178] + error_vector3[179] + error_vector3[180] + error_vector3[181] + error_vector3[182] + error_vector3[183] + error_vector3[184] + error_vector3[185] + error_vector3[186] + error_vector3[187] + error_vector3[188] + error_vector3[189] + error_vector3[190] + error_vector3[191] + error_vector3[192] + error_vector3[193] + error_vector3[194] + error_vector3[195] + error_vector3[196] + error_vector3[197] + error_vector3[198] + error_vector3[199] + error_vector3[200] + error_vector3[201] + error_vector3[202] + error_vector3[203] + error_vector3[204] + error_vector3[205] + error_vector3[206] + error_vector3[207] + error_vector3[208] + error_vector3[209] + error_vector3[210] + error_vector3[211] + error_vector3[212] + error_vector3[213] + error_vector3[214] + error_vector3[215] + error_vector3[216] + error_vector3[217] + error_vector3[218] + error_vector3[219] + error_vector3[220] + error_vector3[221] + error_vector3[222] + error_vector3[223] + error_vector3[224] + error_vector3[225] + error_vector3[226] + error_vector3[227] + error_vector3[228] + error_vector3[229] + error_vector3[230] + error_vector3[231] + error_vector3[232] + error_vector3[233] + error_vector3[234] + error_vector3[235] + error_vector3[236] + error_vector3[237] + error_vector3[238]; 
            errs4 <= error_vector4[0] + error_vector4[1] + error_vector4[2] + error_vector4[3] + error_vector4[4] + error_vector4[5] + error_vector4[6] + error_vector4[7] + error_vector4[8] + error_vector4[9] + error_vector4[10] + error_vector4[11] + error_vector4[12] + error_vector4[13] + error_vector4[14] + error_vector4[15] + error_vector4[16] + error_vector4[17] + error_vector4[18] + error_vector4[19] + error_vector4[20] + error_vector4[21] + error_vector4[22] + error_vector4[23] + error_vector4[24] + error_vector4[25] + error_vector4[26] + error_vector4[27] + error_vector4[28] + error_vector4[29] + error_vector4[30] + error_vector4[31] + error_vector4[32] + error_vector4[33] + error_vector4[34] + error_vector4[35] + error_vector4[36] + error_vector4[37] + error_vector4[38] + error_vector4[39] + error_vector4[40] + error_vector4[41] + error_vector4[42] + error_vector4[43] + error_vector4[44] + error_vector4[45] + error_vector4[46] + error_vector4[47] + error_vector4[48] + error_vector4[49] + error_vector4[50] + error_vector4[51] + error_vector4[52] + error_vector4[53] + error_vector4[54] + error_vector4[55] + error_vector4[56] + error_vector4[57] + error_vector4[58] + error_vector4[59] + error_vector4[60] + error_vector4[61] + error_vector4[62] + error_vector4[63] + error_vector4[64] + error_vector4[65] + error_vector4[66] + error_vector4[67] + error_vector4[68] + error_vector4[69] + error_vector4[70] + error_vector4[71] + error_vector4[72] + error_vector4[73] + error_vector4[74] + error_vector4[75] + error_vector4[76] + error_vector4[77] + error_vector4[78] + error_vector4[79] + error_vector4[80] + error_vector4[81] + error_vector4[82] + error_vector4[83] + error_vector4[84] + error_vector4[85] + error_vector4[86] + error_vector4[87] + error_vector4[88] + error_vector4[89] + error_vector4[90] + error_vector4[91] + error_vector4[92] + error_vector4[93] + error_vector4[94] + error_vector4[95] + error_vector4[96] + error_vector4[97] + error_vector4[98] + error_vector4[99] + error_vector4[100] + error_vector4[101] + error_vector4[102] + error_vector4[103] + error_vector4[104] + error_vector4[105] + error_vector4[106] + error_vector4[107] + error_vector4[108] + error_vector4[109] + error_vector4[110] + error_vector4[111] + error_vector4[112] + error_vector4[113] + error_vector4[114] + error_vector4[115] + error_vector4[116] + error_vector4[117] + error_vector4[118] + error_vector4[119] + error_vector4[120] + error_vector4[121] + error_vector4[122] + error_vector4[123] + error_vector4[124] + error_vector4[125] + error_vector4[126] + error_vector4[127] + error_vector4[128] + error_vector4[129] + error_vector4[130] + error_vector4[131] + error_vector4[132] + error_vector4[133] + error_vector4[134] + error_vector4[135] + error_vector4[136] + error_vector4[137] + error_vector4[138] + error_vector4[139] + error_vector4[140] + error_vector4[141] + error_vector4[142] + error_vector4[143] + error_vector4[144] + error_vector4[145] + error_vector4[146] + error_vector4[147] + error_vector4[148] + error_vector4[149] + error_vector4[150] + error_vector4[151] + error_vector4[152] + error_vector4[153] + error_vector4[154] + error_vector4[155] + error_vector4[156] + error_vector4[157] + error_vector4[158] + error_vector4[159] + error_vector4[160] + error_vector4[161] + error_vector4[162] + error_vector4[163] + error_vector4[164] + error_vector4[165] + error_vector4[166] + error_vector4[167] + error_vector4[168] + error_vector4[169] + error_vector4[170] + error_vector4[171] + error_vector4[172] + error_vector4[173] + error_vector4[174] + error_vector4[175] + error_vector4[176] + error_vector4[177] + error_vector4[178] + error_vector4[179] + error_vector4[180] + error_vector4[181] + error_vector4[182] + error_vector4[183] + error_vector4[184] + error_vector4[185] + error_vector4[186] + error_vector4[187] + error_vector4[188] + error_vector4[189] + error_vector4[190] + error_vector4[191] + error_vector4[192] + error_vector4[193] + error_vector4[194] + error_vector4[195] + error_vector4[196] + error_vector4[197] + error_vector4[198] + error_vector4[199] + error_vector4[200] + error_vector4[201] + error_vector4[202] + error_vector4[203] + error_vector4[204] + error_vector4[205] + error_vector4[206] + error_vector4[207] + error_vector4[208] + error_vector4[209] + error_vector4[210] + error_vector4[211] + error_vector4[212] + error_vector4[213] + error_vector4[214] + error_vector4[215] + error_vector4[216] + error_vector4[217] + error_vector4[218] + error_vector4[219] + error_vector4[220] + error_vector4[221] + error_vector4[222] + error_vector4[223] + error_vector4[224] + error_vector4[225] + error_vector4[226] + error_vector4[227] + error_vector4[228] + error_vector4[229] + error_vector4[230] + error_vector4[231] + error_vector4[232] + error_vector4[233] + error_vector4[234] + error_vector4[235] + error_vector4[236] + error_vector4[237] + error_vector4[238]; 
            errs5 <= error_vector5[0] + error_vector5[1] + error_vector5[2] + error_vector5[3] + error_vector5[4] + error_vector5[5] + error_vector5[6] + error_vector5[7] + error_vector5[8] + error_vector5[9] + error_vector5[10] + error_vector5[11] + error_vector5[12] + error_vector5[13] + error_vector5[14] + error_vector5[15] + error_vector5[16] + error_vector5[17] + error_vector5[18] + error_vector5[19] + error_vector5[20] + error_vector5[21] + error_vector5[22] + error_vector5[23] + error_vector5[24] + error_vector5[25] + error_vector5[26] + error_vector5[27] + error_vector5[28] + error_vector5[29] + error_vector5[30] + error_vector5[31] + error_vector5[32] + error_vector5[33] + error_vector5[34] + error_vector5[35] + error_vector5[36] + error_vector5[37] + error_vector5[38] + error_vector5[39] + error_vector5[40] + error_vector5[41] + error_vector5[42] + error_vector5[43] + error_vector5[44] + error_vector5[45] + error_vector5[46] + error_vector5[47] + error_vector5[48] + error_vector5[49] + error_vector5[50] + error_vector5[51] + error_vector5[52] + error_vector5[53] + error_vector5[54] + error_vector5[55] + error_vector5[56] + error_vector5[57] + error_vector5[58] + error_vector5[59] + error_vector5[60] + error_vector5[61] + error_vector5[62] + error_vector5[63] + error_vector5[64] + error_vector5[65] + error_vector5[66] + error_vector5[67] + error_vector5[68] + error_vector5[69] + error_vector5[70] + error_vector5[71] + error_vector5[72] + error_vector5[73] + error_vector5[74] + error_vector5[75] + error_vector5[76] + error_vector5[77] + error_vector5[78] + error_vector5[79] + error_vector5[80] + error_vector5[81] + error_vector5[82] + error_vector5[83] + error_vector5[84] + error_vector5[85] + error_vector5[86] + error_vector5[87] + error_vector5[88] + error_vector5[89] + error_vector5[90] + error_vector5[91] + error_vector5[92] + error_vector5[93] + error_vector5[94] + error_vector5[95] + error_vector5[96] + error_vector5[97] + error_vector5[98] + error_vector5[99] + error_vector5[100] + error_vector5[101] + error_vector5[102] + error_vector5[103] + error_vector5[104] + error_vector5[105] + error_vector5[106] + error_vector5[107] + error_vector5[108] + error_vector5[109] + error_vector5[110] + error_vector5[111] + error_vector5[112] + error_vector5[113] + error_vector5[114] + error_vector5[115] + error_vector5[116] + error_vector5[117] + error_vector5[118] + error_vector5[119] + error_vector5[120] + error_vector5[121] + error_vector5[122] + error_vector5[123] + error_vector5[124] + error_vector5[125] + error_vector5[126] + error_vector5[127] + error_vector5[128] + error_vector5[129] + error_vector5[130] + error_vector5[131] + error_vector5[132] + error_vector5[133] + error_vector5[134] + error_vector5[135] + error_vector5[136] + error_vector5[137] + error_vector5[138] + error_vector5[139] + error_vector5[140] + error_vector5[141] + error_vector5[142] + error_vector5[143] + error_vector5[144] + error_vector5[145] + error_vector5[146] + error_vector5[147] + error_vector5[148] + error_vector5[149] + error_vector5[150] + error_vector5[151] + error_vector5[152] + error_vector5[153] + error_vector5[154] + error_vector5[155] + error_vector5[156] + error_vector5[157] + error_vector5[158] + error_vector5[159] + error_vector5[160] + error_vector5[161] + error_vector5[162] + error_vector5[163] + error_vector5[164] + error_vector5[165] + error_vector5[166] + error_vector5[167] + error_vector5[168] + error_vector5[169] + error_vector5[170] + error_vector5[171] + error_vector5[172] + error_vector5[173] + error_vector5[174] + error_vector5[175] + error_vector5[176] + error_vector5[177] + error_vector5[178] + error_vector5[179] + error_vector5[180] + error_vector5[181] + error_vector5[182] + error_vector5[183] + error_vector5[184] + error_vector5[185] + error_vector5[186] + error_vector5[187] + error_vector5[188] + error_vector5[189] + error_vector5[190] + error_vector5[191] + error_vector5[192] + error_vector5[193] + error_vector5[194] + error_vector5[195] + error_vector5[196] + error_vector5[197] + error_vector5[198] + error_vector5[199] + error_vector5[200] + error_vector5[201] + error_vector5[202] + error_vector5[203] + error_vector5[204] + error_vector5[205] + error_vector5[206] + error_vector5[207] + error_vector5[208] + error_vector5[209] + error_vector5[210] + error_vector5[211] + error_vector5[212] + error_vector5[213] + error_vector5[214] + error_vector5[215] + error_vector5[216] + error_vector5[217] + error_vector5[218] + error_vector5[219] + error_vector5[220] + error_vector5[221] + error_vector5[222] + error_vector5[223] + error_vector5[224] + error_vector5[225] + error_vector5[226] + error_vector5[227] + error_vector5[228] + error_vector5[229] + error_vector5[230] + error_vector5[231] + error_vector5[232] + error_vector5[233] + error_vector5[234] + error_vector5[235] + error_vector5[236] + error_vector5[237] + error_vector5[238]; 
            errs6 <= error_vector6[0] + error_vector6[1] + error_vector6[2] + error_vector6[3] + error_vector6[4] + error_vector6[5] + error_vector6[6] + error_vector6[7] + error_vector6[8] + error_vector6[9] + error_vector6[10] + error_vector6[11] + error_vector6[12] + error_vector6[13] + error_vector6[14] + error_vector6[15] + error_vector6[16] + error_vector6[17] + error_vector6[18] + error_vector6[19] + error_vector6[20] + error_vector6[21] + error_vector6[22] + error_vector6[23] + error_vector6[24] + error_vector6[25] + error_vector6[26] + error_vector6[27] + error_vector6[28] + error_vector6[29] + error_vector6[30] + error_vector6[31] + error_vector6[32] + error_vector6[33] + error_vector6[34] + error_vector6[35] + error_vector6[36] + error_vector6[37] + error_vector6[38] + error_vector6[39] + error_vector6[40] + error_vector6[41] + error_vector6[42] + error_vector6[43] + error_vector6[44] + error_vector6[45] + error_vector6[46] + error_vector6[47] + error_vector6[48] + error_vector6[49] + error_vector6[50] + error_vector6[51] + error_vector6[52] + error_vector6[53] + error_vector6[54] + error_vector6[55] + error_vector6[56] + error_vector6[57] + error_vector6[58] + error_vector6[59] + error_vector6[60] + error_vector6[61] + error_vector6[62] + error_vector6[63] + error_vector6[64] + error_vector6[65] + error_vector6[66] + error_vector6[67] + error_vector6[68] + error_vector6[69] + error_vector6[70] + error_vector6[71] + error_vector6[72] + error_vector6[73] + error_vector6[74] + error_vector6[75] + error_vector6[76] + error_vector6[77] + error_vector6[78] + error_vector6[79] + error_vector6[80] + error_vector6[81] + error_vector6[82] + error_vector6[83] + error_vector6[84] + error_vector6[85] + error_vector6[86] + error_vector6[87] + error_vector6[88] + error_vector6[89] + error_vector6[90] + error_vector6[91] + error_vector6[92] + error_vector6[93] + error_vector6[94] + error_vector6[95] + error_vector6[96] + error_vector6[97] + error_vector6[98] + error_vector6[99] + error_vector6[100] + error_vector6[101] + error_vector6[102] + error_vector6[103] + error_vector6[104] + error_vector6[105] + error_vector6[106] + error_vector6[107] + error_vector6[108] + error_vector6[109] + error_vector6[110] + error_vector6[111] + error_vector6[112] + error_vector6[113] + error_vector6[114] + error_vector6[115] + error_vector6[116] + error_vector6[117] + error_vector6[118] + error_vector6[119] + error_vector6[120] + error_vector6[121] + error_vector6[122] + error_vector6[123] + error_vector6[124] + error_vector6[125] + error_vector6[126] + error_vector6[127] + error_vector6[128] + error_vector6[129] + error_vector6[130] + error_vector6[131] + error_vector6[132] + error_vector6[133] + error_vector6[134] + error_vector6[135] + error_vector6[136] + error_vector6[137] + error_vector6[138] + error_vector6[139] + error_vector6[140] + error_vector6[141] + error_vector6[142] + error_vector6[143] + error_vector6[144] + error_vector6[145] + error_vector6[146] + error_vector6[147] + error_vector6[148] + error_vector6[149] + error_vector6[150] + error_vector6[151] + error_vector6[152] + error_vector6[153] + error_vector6[154] + error_vector6[155] + error_vector6[156] + error_vector6[157] + error_vector6[158] + error_vector6[159] + error_vector6[160] + error_vector6[161] + error_vector6[162] + error_vector6[163] + error_vector6[164] + error_vector6[165] + error_vector6[166] + error_vector6[167] + error_vector6[168] + error_vector6[169] + error_vector6[170] + error_vector6[171] + error_vector6[172] + error_vector6[173] + error_vector6[174] + error_vector6[175] + error_vector6[176] + error_vector6[177] + error_vector6[178] + error_vector6[179] + error_vector6[180] + error_vector6[181] + error_vector6[182] + error_vector6[183] + error_vector6[184] + error_vector6[185] + error_vector6[186] + error_vector6[187] + error_vector6[188] + error_vector6[189] + error_vector6[190] + error_vector6[191] + error_vector6[192] + error_vector6[193] + error_vector6[194] + error_vector6[195] + error_vector6[196] + error_vector6[197] + error_vector6[198] + error_vector6[199] + error_vector6[200] + error_vector6[201] + error_vector6[202] + error_vector6[203] + error_vector6[204] + error_vector6[205] + error_vector6[206] + error_vector6[207] + error_vector6[208] + error_vector6[209] + error_vector6[210] + error_vector6[211] + error_vector6[212] + error_vector6[213] + error_vector6[214] + error_vector6[215] + error_vector6[216] + error_vector6[217] + error_vector6[218] + error_vector6[219] + error_vector6[220] + error_vector6[221] + error_vector6[222] + error_vector6[223] + error_vector6[224] + error_vector6[225] + error_vector6[226] + error_vector6[227] + error_vector6[228] + error_vector6[229] + error_vector6[230] + error_vector6[231] + error_vector6[232] + error_vector6[233] + error_vector6[234] + error_vector6[235] + error_vector6[236] + error_vector6[237] + error_vector6[238]; 
            errs7 <= error_vector7[0] + error_vector7[1] + error_vector7[2] + error_vector7[3] + error_vector7[4] + error_vector7[5] + error_vector7[6] + error_vector7[7] + error_vector7[8] + error_vector7[9] + error_vector7[10] + error_vector7[11] + error_vector7[12] + error_vector7[13] + error_vector7[14] + error_vector7[15] + error_vector7[16] + error_vector7[17] + error_vector7[18] + error_vector7[19] + error_vector7[20] + error_vector7[21] + error_vector7[22] + error_vector7[23] + error_vector7[24] + error_vector7[25] + error_vector7[26] + error_vector7[27] + error_vector7[28] + error_vector7[29] + error_vector7[30] + error_vector7[31] + error_vector7[32] + error_vector7[33] + error_vector7[34] + error_vector7[35] + error_vector7[36] + error_vector7[37] + error_vector7[38] + error_vector7[39] + error_vector7[40] + error_vector7[41] + error_vector7[42] + error_vector7[43] + error_vector7[44] + error_vector7[45] + error_vector7[46] + error_vector7[47] + error_vector7[48] + error_vector7[49] + error_vector7[50] + error_vector7[51] + error_vector7[52] + error_vector7[53] + error_vector7[54] + error_vector7[55] + error_vector7[56] + error_vector7[57] + error_vector7[58] + error_vector7[59] + error_vector7[60] + error_vector7[61] + error_vector7[62] + error_vector7[63] + error_vector7[64] + error_vector7[65] + error_vector7[66] + error_vector7[67] + error_vector7[68] + error_vector7[69] + error_vector7[70] + error_vector7[71] + error_vector7[72] + error_vector7[73] + error_vector7[74] + error_vector7[75] + error_vector7[76] + error_vector7[77] + error_vector7[78] + error_vector7[79] + error_vector7[80] + error_vector7[81] + error_vector7[82] + error_vector7[83] + error_vector7[84] + error_vector7[85] + error_vector7[86] + error_vector7[87] + error_vector7[88] + error_vector7[89] + error_vector7[90] + error_vector7[91] + error_vector7[92] + error_vector7[93] + error_vector7[94] + error_vector7[95] + error_vector7[96] + error_vector7[97] + error_vector7[98] + error_vector7[99] + error_vector7[100] + error_vector7[101] + error_vector7[102] + error_vector7[103] + error_vector7[104] + error_vector7[105] + error_vector7[106] + error_vector7[107] + error_vector7[108] + error_vector7[109] + error_vector7[110] + error_vector7[111] + error_vector7[112] + error_vector7[113] + error_vector7[114] + error_vector7[115] + error_vector7[116] + error_vector7[117] + error_vector7[118] + error_vector7[119] + error_vector7[120] + error_vector7[121] + error_vector7[122] + error_vector7[123] + error_vector7[124] + error_vector7[125] + error_vector7[126] + error_vector7[127] + error_vector7[128] + error_vector7[129] + error_vector7[130] + error_vector7[131] + error_vector7[132] + error_vector7[133] + error_vector7[134] + error_vector7[135] + error_vector7[136] + error_vector7[137] + error_vector7[138] + error_vector7[139] + error_vector7[140] + error_vector7[141] + error_vector7[142] + error_vector7[143] + error_vector7[144] + error_vector7[145] + error_vector7[146] + error_vector7[147] + error_vector7[148] + error_vector7[149] + error_vector7[150] + error_vector7[151] + error_vector7[152] + error_vector7[153] + error_vector7[154] + error_vector7[155] + error_vector7[156] + error_vector7[157] + error_vector7[158] + error_vector7[159] + error_vector7[160] + error_vector7[161] + error_vector7[162] + error_vector7[163] + error_vector7[164] + error_vector7[165] + error_vector7[166] + error_vector7[167] + error_vector7[168] + error_vector7[169] + error_vector7[170] + error_vector7[171] + error_vector7[172] + error_vector7[173] + error_vector7[174] + error_vector7[175] + error_vector7[176] + error_vector7[177] + error_vector7[178] + error_vector7[179] + error_vector7[180] + error_vector7[181] + error_vector7[182] + error_vector7[183] + error_vector7[184] + error_vector7[185] + error_vector7[186] + error_vector7[187] + error_vector7[188] + error_vector7[189] + error_vector7[190] + error_vector7[191] + error_vector7[192] + error_vector7[193] + error_vector7[194] + error_vector7[195] + error_vector7[196] + error_vector7[197] + error_vector7[198] + error_vector7[199] + error_vector7[200] + error_vector7[201] + error_vector7[202] + error_vector7[203] + error_vector7[204] + error_vector7[205] + error_vector7[206] + error_vector7[207] + error_vector7[208] + error_vector7[209] + error_vector7[210] + error_vector7[211] + error_vector7[212] + error_vector7[213] + error_vector7[214] + error_vector7[215] + error_vector7[216] + error_vector7[217] + error_vector7[218] + error_vector7[219] + error_vector7[220] + error_vector7[221] + error_vector7[222] + error_vector7[223] + error_vector7[224] + error_vector7[225] + error_vector7[226] + error_vector7[227] + error_vector7[228] + error_vector7[229] + error_vector7[230] + error_vector7[231] + error_vector7[232] + error_vector7[233] + error_vector7[234] + error_vector7[235] + error_vector7[236] + error_vector7[237] + error_vector7[238]; 
            errs8 <= error_vector8[0] + error_vector8[1] + error_vector8[2] + error_vector8[3] + error_vector8[4] + error_vector8[5] + error_vector8[6] + error_vector8[7] + error_vector8[8] + error_vector8[9] + error_vector8[10] + error_vector8[11] + error_vector8[12] + error_vector8[13] + error_vector8[14] + error_vector8[15] + error_vector8[16] + error_vector8[17] + error_vector8[18] + error_vector8[19] + error_vector8[20] + error_vector8[21] + error_vector8[22] + error_vector8[23] + error_vector8[24] + error_vector8[25] + error_vector8[26] + error_vector8[27] + error_vector8[28] + error_vector8[29] + error_vector8[30] + error_vector8[31] + error_vector8[32] + error_vector8[33] + error_vector8[34] + error_vector8[35] + error_vector8[36] + error_vector8[37] + error_vector8[38] + error_vector8[39] + error_vector8[40] + error_vector8[41] + error_vector8[42] + error_vector8[43] + error_vector8[44] + error_vector8[45] + error_vector8[46] + error_vector8[47] + error_vector8[48] + error_vector8[49] + error_vector8[50] + error_vector8[51] + error_vector8[52] + error_vector8[53] + error_vector8[54] + error_vector8[55] + error_vector8[56] + error_vector8[57] + error_vector8[58] + error_vector8[59] + error_vector8[60] + error_vector8[61] + error_vector8[62] + error_vector8[63] + error_vector8[64] + error_vector8[65] + error_vector8[66] + error_vector8[67] + error_vector8[68] + error_vector8[69] + error_vector8[70] + error_vector8[71] + error_vector8[72] + error_vector8[73] + error_vector8[74] + error_vector8[75] + error_vector8[76] + error_vector8[77] + error_vector8[78] + error_vector8[79] + error_vector8[80] + error_vector8[81] + error_vector8[82] + error_vector8[83] + error_vector8[84] + error_vector8[85] + error_vector8[86] + error_vector8[87] + error_vector8[88] + error_vector8[89] + error_vector8[90] + error_vector8[91] + error_vector8[92] + error_vector8[93] + error_vector8[94] + error_vector8[95] + error_vector8[96] + error_vector8[97] + error_vector8[98] + error_vector8[99] + error_vector8[100] + error_vector8[101] + error_vector8[102] + error_vector8[103] + error_vector8[104] + error_vector8[105] + error_vector8[106] + error_vector8[107] + error_vector8[108] + error_vector8[109] + error_vector8[110] + error_vector8[111] + error_vector8[112] + error_vector8[113] + error_vector8[114] + error_vector8[115] + error_vector8[116] + error_vector8[117] + error_vector8[118] + error_vector8[119] + error_vector8[120] + error_vector8[121] + error_vector8[122] + error_vector8[123] + error_vector8[124] + error_vector8[125] + error_vector8[126] + error_vector8[127] + error_vector8[128] + error_vector8[129] + error_vector8[130] + error_vector8[131] + error_vector8[132] + error_vector8[133] + error_vector8[134] + error_vector8[135] + error_vector8[136] + error_vector8[137] + error_vector8[138] + error_vector8[139] + error_vector8[140] + error_vector8[141] + error_vector8[142] + error_vector8[143] + error_vector8[144] + error_vector8[145] + error_vector8[146] + error_vector8[147] + error_vector8[148] + error_vector8[149] + error_vector8[150] + error_vector8[151] + error_vector8[152] + error_vector8[153] + error_vector8[154] + error_vector8[155] + error_vector8[156] + error_vector8[157] + error_vector8[158] + error_vector8[159] + error_vector8[160] + error_vector8[161] + error_vector8[162] + error_vector8[163] + error_vector8[164] + error_vector8[165] + error_vector8[166] + error_vector8[167] + error_vector8[168] + error_vector8[169] + error_vector8[170] + error_vector8[171] + error_vector8[172] + error_vector8[173] + error_vector8[174] + error_vector8[175] + error_vector8[176] + error_vector8[177] + error_vector8[178] + error_vector8[179] + error_vector8[180] + error_vector8[181] + error_vector8[182] + error_vector8[183] + error_vector8[184] + error_vector8[185] + error_vector8[186] + error_vector8[187] + error_vector8[188] + error_vector8[189] + error_vector8[190] + error_vector8[191] + error_vector8[192] + error_vector8[193] + error_vector8[194] + error_vector8[195] + error_vector8[196] + error_vector8[197] + error_vector8[198] + error_vector8[199] + error_vector8[200] + error_vector8[201] + error_vector8[202] + error_vector8[203] + error_vector8[204] + error_vector8[205] + error_vector8[206] + error_vector8[207] + error_vector8[208] + error_vector8[209] + error_vector8[210] + error_vector8[211] + error_vector8[212] + error_vector8[213] + error_vector8[214] + error_vector8[215] + error_vector8[216] + error_vector8[217] + error_vector8[218] + error_vector8[219] + error_vector8[220] + error_vector8[221] + error_vector8[222] + error_vector8[223] + error_vector8[224] + error_vector8[225] + error_vector8[226] + error_vector8[227] + error_vector8[228] + error_vector8[229] + error_vector8[230] + error_vector8[231] + error_vector8[232] + error_vector8[233] + error_vector8[234] + error_vector8[235] + error_vector8[236] + error_vector8[237] + error_vector8[238]; 
            errs9 <= error_vector9[0] + error_vector9[1] + error_vector9[2] + error_vector9[3] + error_vector9[4] + error_vector9[5] + error_vector9[6] + error_vector9[7] + error_vector9[8] + error_vector9[9] + error_vector9[10] + error_vector9[11] + error_vector9[12] + error_vector9[13] + error_vector9[14] + error_vector9[15] + error_vector9[16] + error_vector9[17] + error_vector9[18] + error_vector9[19] + error_vector9[20] + error_vector9[21] + error_vector9[22] + error_vector9[23] + error_vector9[24] + error_vector9[25] + error_vector9[26] + error_vector9[27] + error_vector9[28] + error_vector9[29] + error_vector9[30] + error_vector9[31] + error_vector9[32] + error_vector9[33] + error_vector9[34] + error_vector9[35] + error_vector9[36] + error_vector9[37] + error_vector9[38] + error_vector9[39] + error_vector9[40] + error_vector9[41] + error_vector9[42] + error_vector9[43] + error_vector9[44] + error_vector9[45] + error_vector9[46] + error_vector9[47] + error_vector9[48] + error_vector9[49] + error_vector9[50] + error_vector9[51] + error_vector9[52] + error_vector9[53] + error_vector9[54] + error_vector9[55] + error_vector9[56] + error_vector9[57] + error_vector9[58] + error_vector9[59] + error_vector9[60] + error_vector9[61] + error_vector9[62] + error_vector9[63] + error_vector9[64] + error_vector9[65] + error_vector9[66] + error_vector9[67] + error_vector9[68] + error_vector9[69] + error_vector9[70] + error_vector9[71] + error_vector9[72] + error_vector9[73] + error_vector9[74] + error_vector9[75] + error_vector9[76] + error_vector9[77] + error_vector9[78] + error_vector9[79] + error_vector9[80] + error_vector9[81] + error_vector9[82] + error_vector9[83] + error_vector9[84] + error_vector9[85] + error_vector9[86] + error_vector9[87] + error_vector9[88] + error_vector9[89] + error_vector9[90] + error_vector9[91] + error_vector9[92] + error_vector9[93] + error_vector9[94] + error_vector9[95] + error_vector9[96] + error_vector9[97] + error_vector9[98] + error_vector9[99] + error_vector9[100] + error_vector9[101] + error_vector9[102] + error_vector9[103] + error_vector9[104] + error_vector9[105] + error_vector9[106] + error_vector9[107] + error_vector9[108] + error_vector9[109] + error_vector9[110] + error_vector9[111] + error_vector9[112] + error_vector9[113] + error_vector9[114] + error_vector9[115] + error_vector9[116] + error_vector9[117] + error_vector9[118] + error_vector9[119] + error_vector9[120] + error_vector9[121] + error_vector9[122] + error_vector9[123] + error_vector9[124] + error_vector9[125] + error_vector9[126] + error_vector9[127] + error_vector9[128] + error_vector9[129] + error_vector9[130] + error_vector9[131] + error_vector9[132] + error_vector9[133] + error_vector9[134] + error_vector9[135] + error_vector9[136] + error_vector9[137] + error_vector9[138] + error_vector9[139] + error_vector9[140] + error_vector9[141] + error_vector9[142] + error_vector9[143] + error_vector9[144] + error_vector9[145] + error_vector9[146] + error_vector9[147] + error_vector9[148] + error_vector9[149] + error_vector9[150] + error_vector9[151] + error_vector9[152] + error_vector9[153] + error_vector9[154] + error_vector9[155] + error_vector9[156] + error_vector9[157] + error_vector9[158] + error_vector9[159] + error_vector9[160] + error_vector9[161] + error_vector9[162] + error_vector9[163] + error_vector9[164] + error_vector9[165] + error_vector9[166] + error_vector9[167] + error_vector9[168] + error_vector9[169] + error_vector9[170] + error_vector9[171] + error_vector9[172] + error_vector9[173] + error_vector9[174] + error_vector9[175] + error_vector9[176] + error_vector9[177] + error_vector9[178] + error_vector9[179] + error_vector9[180] + error_vector9[181] + error_vector9[182] + error_vector9[183] + error_vector9[184] + error_vector9[185] + error_vector9[186] + error_vector9[187] + error_vector9[188] + error_vector9[189] + error_vector9[190] + error_vector9[191] + error_vector9[192] + error_vector9[193] + error_vector9[194] + error_vector9[195] + error_vector9[196] + error_vector9[197] + error_vector9[198] + error_vector9[199] + error_vector9[200] + error_vector9[201] + error_vector9[202] + error_vector9[203] + error_vector9[204] + error_vector9[205] + error_vector9[206] + error_vector9[207] + error_vector9[208] + error_vector9[209] + error_vector9[210] + error_vector9[211] + error_vector9[212] + error_vector9[213] + error_vector9[214] + error_vector9[215] + error_vector9[216] + error_vector9[217] + error_vector9[218] + error_vector9[219] + error_vector9[220] + error_vector9[221] + error_vector9[222] + error_vector9[223] + error_vector9[224] + error_vector9[225] + error_vector9[226] + error_vector9[227] + error_vector9[228] + error_vector9[229] + error_vector9[230] + error_vector9[231] + error_vector9[232] + error_vector9[233] + error_vector9[234] + error_vector9[235] + error_vector9[236] + error_vector9[237] + error_vector9[238]; 
            errs10 <= error_vector10[0] + error_vector10[1] + error_vector10[2] + error_vector10[3] + error_vector10[4] + error_vector10[5] + error_vector10[6] + error_vector10[7] + error_vector10[8] + error_vector10[9] + error_vector10[10] + error_vector10[11] + error_vector10[12] + error_vector10[13] + error_vector10[14] + error_vector10[15] + error_vector10[16] + error_vector10[17] + error_vector10[18] + error_vector10[19] + error_vector10[20] + error_vector10[21] + error_vector10[22] + error_vector10[23] + error_vector10[24] + error_vector10[25] + error_vector10[26] + error_vector10[27] + error_vector10[28] + error_vector10[29] + error_vector10[30] + error_vector10[31] + error_vector10[32] + error_vector10[33] + error_vector10[34] + error_vector10[35] + error_vector10[36] + error_vector10[37] + error_vector10[38] + error_vector10[39] + error_vector10[40] + error_vector10[41] + error_vector10[42] + error_vector10[43] + error_vector10[44] + error_vector10[45] + error_vector10[46] + error_vector10[47] + error_vector10[48] + error_vector10[49] + error_vector10[50] + error_vector10[51] + error_vector10[52] + error_vector10[53] + error_vector10[54] + error_vector10[55] + error_vector10[56] + error_vector10[57] + error_vector10[58] + error_vector10[59] + error_vector10[60] + error_vector10[61] + error_vector10[62] + error_vector10[63] + error_vector10[64] + error_vector10[65] + error_vector10[66] + error_vector10[67] + error_vector10[68] + error_vector10[69] + error_vector10[70] + error_vector10[71] + error_vector10[72] + error_vector10[73] + error_vector10[74] + error_vector10[75] + error_vector10[76] + error_vector10[77] + error_vector10[78] + error_vector10[79] + error_vector10[80] + error_vector10[81] + error_vector10[82] + error_vector10[83] + error_vector10[84] + error_vector10[85] + error_vector10[86] + error_vector10[87] + error_vector10[88] + error_vector10[89] + error_vector10[90] + error_vector10[91] + error_vector10[92] + error_vector10[93] + error_vector10[94] + error_vector10[95] + error_vector10[96] + error_vector10[97] + error_vector10[98] + error_vector10[99] + error_vector10[100] + error_vector10[101] + error_vector10[102] + error_vector10[103] + error_vector10[104] + error_vector10[105] + error_vector10[106] + error_vector10[107] + error_vector10[108] + error_vector10[109] + error_vector10[110] + error_vector10[111] + error_vector10[112] + error_vector10[113] + error_vector10[114] + error_vector10[115] + error_vector10[116] + error_vector10[117] + error_vector10[118] + error_vector10[119] + error_vector10[120] + error_vector10[121] + error_vector10[122] + error_vector10[123] + error_vector10[124] + error_vector10[125] + error_vector10[126] + error_vector10[127] + error_vector10[128] + error_vector10[129] + error_vector10[130] + error_vector10[131] + error_vector10[132] + error_vector10[133] + error_vector10[134] + error_vector10[135] + error_vector10[136] + error_vector10[137] + error_vector10[138] + error_vector10[139] + error_vector10[140] + error_vector10[141] + error_vector10[142] + error_vector10[143] + error_vector10[144] + error_vector10[145] + error_vector10[146] + error_vector10[147] + error_vector10[148] + error_vector10[149] + error_vector10[150] + error_vector10[151] + error_vector10[152] + error_vector10[153] + error_vector10[154] + error_vector10[155] + error_vector10[156] + error_vector10[157] + error_vector10[158] + error_vector10[159] + error_vector10[160] + error_vector10[161] + error_vector10[162] + error_vector10[163] + error_vector10[164] + error_vector10[165] + error_vector10[166] + error_vector10[167] + error_vector10[168] + error_vector10[169] + error_vector10[170] + error_vector10[171] + error_vector10[172] + error_vector10[173] + error_vector10[174] + error_vector10[175] + error_vector10[176] + error_vector10[177] + error_vector10[178] + error_vector10[179] + error_vector10[180] + error_vector10[181] + error_vector10[182] + error_vector10[183] + error_vector10[184] + error_vector10[185] + error_vector10[186] + error_vector10[187] + error_vector10[188] + error_vector10[189] + error_vector10[190] + error_vector10[191] + error_vector10[192] + error_vector10[193] + error_vector10[194] + error_vector10[195] + error_vector10[196] + error_vector10[197] + error_vector10[198] + error_vector10[199] + error_vector10[200] + error_vector10[201] + error_vector10[202] + error_vector10[203] + error_vector10[204] + error_vector10[205] + error_vector10[206] + error_vector10[207] + error_vector10[208] + error_vector10[209] + error_vector10[210] + error_vector10[211] + error_vector10[212] + error_vector10[213] + error_vector10[214] + error_vector10[215] + error_vector10[216] + error_vector10[217] + error_vector10[218] + error_vector10[219] + error_vector10[220] + error_vector10[221] + error_vector10[222] + error_vector10[223] + error_vector10[224] + error_vector10[225] + error_vector10[226] + error_vector10[227] + error_vector10[228] + error_vector10[229] + error_vector10[230] + error_vector10[231] + error_vector10[232] + error_vector10[233] + error_vector10[234] + error_vector10[235] + error_vector10[236] + error_vector10[237] + error_vector10[238]; 
            errs11 <= error_vector11[0] + error_vector11[1] + error_vector11[2] + error_vector11[3] + error_vector11[4] + error_vector11[5] + error_vector11[6] + error_vector11[7] + error_vector11[8] + error_vector11[9] + error_vector11[10] + error_vector11[11] + error_vector11[12] + error_vector11[13] + error_vector11[14] + error_vector11[15] + error_vector11[16] + error_vector11[17] + error_vector11[18] + error_vector11[19] + error_vector11[20] + error_vector11[21] + error_vector11[22] + error_vector11[23] + error_vector11[24] + error_vector11[25] + error_vector11[26] + error_vector11[27] + error_vector11[28] + error_vector11[29] + error_vector11[30] + error_vector11[31] + error_vector11[32] + error_vector11[33] + error_vector11[34] + error_vector11[35] + error_vector11[36] + error_vector11[37] + error_vector11[38] + error_vector11[39] + error_vector11[40] + error_vector11[41] + error_vector11[42] + error_vector11[43] + error_vector11[44] + error_vector11[45] + error_vector11[46] + error_vector11[47] + error_vector11[48] + error_vector11[49] + error_vector11[50] + error_vector11[51] + error_vector11[52] + error_vector11[53] + error_vector11[54] + error_vector11[55] + error_vector11[56] + error_vector11[57] + error_vector11[58] + error_vector11[59] + error_vector11[60] + error_vector11[61] + error_vector11[62] + error_vector11[63] + error_vector11[64] + error_vector11[65] + error_vector11[66] + error_vector11[67] + error_vector11[68] + error_vector11[69] + error_vector11[70] + error_vector11[71] + error_vector11[72] + error_vector11[73] + error_vector11[74] + error_vector11[75] + error_vector11[76] + error_vector11[77] + error_vector11[78] + error_vector11[79] + error_vector11[80] + error_vector11[81] + error_vector11[82] + error_vector11[83] + error_vector11[84] + error_vector11[85] + error_vector11[86] + error_vector11[87] + error_vector11[88] + error_vector11[89] + error_vector11[90] + error_vector11[91] + error_vector11[92] + error_vector11[93] + error_vector11[94] + error_vector11[95] + error_vector11[96] + error_vector11[97] + error_vector11[98] + error_vector11[99] + error_vector11[100] + error_vector11[101] + error_vector11[102] + error_vector11[103] + error_vector11[104] + error_vector11[105] + error_vector11[106] + error_vector11[107] + error_vector11[108] + error_vector11[109] + error_vector11[110] + error_vector11[111] + error_vector11[112] + error_vector11[113] + error_vector11[114] + error_vector11[115] + error_vector11[116] + error_vector11[117] + error_vector11[118] + error_vector11[119] + error_vector11[120] + error_vector11[121] + error_vector11[122] + error_vector11[123] + error_vector11[124] + error_vector11[125] + error_vector11[126] + error_vector11[127] + error_vector11[128] + error_vector11[129] + error_vector11[130] + error_vector11[131] + error_vector11[132] + error_vector11[133] + error_vector11[134] + error_vector11[135] + error_vector11[136] + error_vector11[137] + error_vector11[138] + error_vector11[139] + error_vector11[140] + error_vector11[141] + error_vector11[142] + error_vector11[143] + error_vector11[144] + error_vector11[145] + error_vector11[146] + error_vector11[147] + error_vector11[148] + error_vector11[149] + error_vector11[150] + error_vector11[151] + error_vector11[152] + error_vector11[153] + error_vector11[154] + error_vector11[155] + error_vector11[156] + error_vector11[157] + error_vector11[158] + error_vector11[159] + error_vector11[160] + error_vector11[161] + error_vector11[162] + error_vector11[163] + error_vector11[164] + error_vector11[165] + error_vector11[166] + error_vector11[167] + error_vector11[168] + error_vector11[169] + error_vector11[170] + error_vector11[171] + error_vector11[172] + error_vector11[173] + error_vector11[174] + error_vector11[175] + error_vector11[176] + error_vector11[177] + error_vector11[178] + error_vector11[179] + error_vector11[180] + error_vector11[181] + error_vector11[182] + error_vector11[183] + error_vector11[184] + error_vector11[185] + error_vector11[186] + error_vector11[187] + error_vector11[188] + error_vector11[189] + error_vector11[190] + error_vector11[191] + error_vector11[192] + error_vector11[193] + error_vector11[194] + error_vector11[195] + error_vector11[196] + error_vector11[197] + error_vector11[198] + error_vector11[199] + error_vector11[200] + error_vector11[201] + error_vector11[202] + error_vector11[203] + error_vector11[204] + error_vector11[205] + error_vector11[206] + error_vector11[207] + error_vector11[208] + error_vector11[209] + error_vector11[210] + error_vector11[211] + error_vector11[212] + error_vector11[213] + error_vector11[214] + error_vector11[215] + error_vector11[216] + error_vector11[217] + error_vector11[218] + error_vector11[219] + error_vector11[220] + error_vector11[221] + error_vector11[222] + error_vector11[223] + error_vector11[224] + error_vector11[225] + error_vector11[226] + error_vector11[227] + error_vector11[228] + error_vector11[229] + error_vector11[230] + error_vector11[231] + error_vector11[232] + error_vector11[233] + error_vector11[234] + error_vector11[235] + error_vector11[236] + error_vector11[237] + error_vector11[238]; 
            errs12 <= error_vector12[0] + error_vector12[1] + error_vector12[2] + error_vector12[3] + error_vector12[4] + error_vector12[5] + error_vector12[6] + error_vector12[7] + error_vector12[8] + error_vector12[9] + error_vector12[10] + error_vector12[11] + error_vector12[12] + error_vector12[13] + error_vector12[14] + error_vector12[15] + error_vector12[16] + error_vector12[17] + error_vector12[18] + error_vector12[19] + error_vector12[20] + error_vector12[21] + error_vector12[22] + error_vector12[23] + error_vector12[24] + error_vector12[25] + error_vector12[26] + error_vector12[27] + error_vector12[28] + error_vector12[29] + error_vector12[30] + error_vector12[31] + error_vector12[32] + error_vector12[33] + error_vector12[34] + error_vector12[35] + error_vector12[36] + error_vector12[37] + error_vector12[38] + error_vector12[39] + error_vector12[40] + error_vector12[41] + error_vector12[42] + error_vector12[43] + error_vector12[44] + error_vector12[45] + error_vector12[46] + error_vector12[47] + error_vector12[48] + error_vector12[49] + error_vector12[50] + error_vector12[51] + error_vector12[52] + error_vector12[53] + error_vector12[54] + error_vector12[55] + error_vector12[56] + error_vector12[57] + error_vector12[58] + error_vector12[59] + error_vector12[60] + error_vector12[61] + error_vector12[62] + error_vector12[63] + error_vector12[64] + error_vector12[65] + error_vector12[66] + error_vector12[67] + error_vector12[68] + error_vector12[69] + error_vector12[70] + error_vector12[71] + error_vector12[72] + error_vector12[73] + error_vector12[74] + error_vector12[75] + error_vector12[76] + error_vector12[77] + error_vector12[78] + error_vector12[79] + error_vector12[80] + error_vector12[81] + error_vector12[82] + error_vector12[83] + error_vector12[84] + error_vector12[85] + error_vector12[86] + error_vector12[87] + error_vector12[88] + error_vector12[89] + error_vector12[90] + error_vector12[91] + error_vector12[92] + error_vector12[93] + error_vector12[94] + error_vector12[95] + error_vector12[96] + error_vector12[97] + error_vector12[98] + error_vector12[99] + error_vector12[100] + error_vector12[101] + error_vector12[102] + error_vector12[103] + error_vector12[104] + error_vector12[105] + error_vector12[106] + error_vector12[107] + error_vector12[108] + error_vector12[109] + error_vector12[110] + error_vector12[111] + error_vector12[112] + error_vector12[113] + error_vector12[114] + error_vector12[115] + error_vector12[116] + error_vector12[117] + error_vector12[118] + error_vector12[119] + error_vector12[120] + error_vector12[121] + error_vector12[122] + error_vector12[123] + error_vector12[124] + error_vector12[125] + error_vector12[126] + error_vector12[127] + error_vector12[128] + error_vector12[129] + error_vector12[130] + error_vector12[131] + error_vector12[132] + error_vector12[133] + error_vector12[134] + error_vector12[135] + error_vector12[136] + error_vector12[137] + error_vector12[138] + error_vector12[139] + error_vector12[140] + error_vector12[141] + error_vector12[142] + error_vector12[143] + error_vector12[144] + error_vector12[145] + error_vector12[146] + error_vector12[147] + error_vector12[148] + error_vector12[149] + error_vector12[150] + error_vector12[151] + error_vector12[152] + error_vector12[153] + error_vector12[154] + error_vector12[155] + error_vector12[156] + error_vector12[157] + error_vector12[158] + error_vector12[159] + error_vector12[160] + error_vector12[161] + error_vector12[162] + error_vector12[163] + error_vector12[164] + error_vector12[165] + error_vector12[166] + error_vector12[167] + error_vector12[168] + error_vector12[169] + error_vector12[170] + error_vector12[171] + error_vector12[172] + error_vector12[173] + error_vector12[174] + error_vector12[175] + error_vector12[176] + error_vector12[177] + error_vector12[178] + error_vector12[179] + error_vector12[180] + error_vector12[181] + error_vector12[182] + error_vector12[183] + error_vector12[184] + error_vector12[185] + error_vector12[186] + error_vector12[187] + error_vector12[188] + error_vector12[189] + error_vector12[190] + error_vector12[191] + error_vector12[192] + error_vector12[193] + error_vector12[194] + error_vector12[195] + error_vector12[196] + error_vector12[197] + error_vector12[198] + error_vector12[199] + error_vector12[200] + error_vector12[201] + error_vector12[202] + error_vector12[203] + error_vector12[204] + error_vector12[205] + error_vector12[206] + error_vector12[207] + error_vector12[208] + error_vector12[209] + error_vector12[210] + error_vector12[211] + error_vector12[212] + error_vector12[213] + error_vector12[214] + error_vector12[215] + error_vector12[216] + error_vector12[217] + error_vector12[218] + error_vector12[219] + error_vector12[220] + error_vector12[221] + error_vector12[222] + error_vector12[223] + error_vector12[224] + error_vector12[225] + error_vector12[226] + error_vector12[227] + error_vector12[228] + error_vector12[229] + error_vector12[230] + error_vector12[231] + error_vector12[232] + error_vector12[233] + error_vector12[234] + error_vector12[235] + error_vector12[236] + error_vector12[237] + error_vector12[238]; 
            errs13 <= error_vector13[0] + error_vector13[1] + error_vector13[2] + error_vector13[3] + error_vector13[4] + error_vector13[5] + error_vector13[6] + error_vector13[7] + error_vector13[8] + error_vector13[9] + error_vector13[10] + error_vector13[11] + error_vector13[12] + error_vector13[13] + error_vector13[14] + error_vector13[15] + error_vector13[16] + error_vector13[17] + error_vector13[18] + error_vector13[19] + error_vector13[20] + error_vector13[21] + error_vector13[22] + error_vector13[23] + error_vector13[24] + error_vector13[25] + error_vector13[26] + error_vector13[27] + error_vector13[28] + error_vector13[29] + error_vector13[30] + error_vector13[31] + error_vector13[32] + error_vector13[33] + error_vector13[34] + error_vector13[35] + error_vector13[36] + error_vector13[37] + error_vector13[38] + error_vector13[39] + error_vector13[40] + error_vector13[41] + error_vector13[42] + error_vector13[43] + error_vector13[44] + error_vector13[45] + error_vector13[46] + error_vector13[47] + error_vector13[48] + error_vector13[49] + error_vector13[50] + error_vector13[51] + error_vector13[52] + error_vector13[53] + error_vector13[54] + error_vector13[55] + error_vector13[56] + error_vector13[57] + error_vector13[58] + error_vector13[59] + error_vector13[60] + error_vector13[61] + error_vector13[62] + error_vector13[63] + error_vector13[64] + error_vector13[65] + error_vector13[66] + error_vector13[67] + error_vector13[68] + error_vector13[69] + error_vector13[70] + error_vector13[71] + error_vector13[72] + error_vector13[73] + error_vector13[74] + error_vector13[75] + error_vector13[76] + error_vector13[77] + error_vector13[78] + error_vector13[79] + error_vector13[80] + error_vector13[81] + error_vector13[82] + error_vector13[83] + error_vector13[84] + error_vector13[85] + error_vector13[86] + error_vector13[87] + error_vector13[88] + error_vector13[89] + error_vector13[90] + error_vector13[91] + error_vector13[92] + error_vector13[93] + error_vector13[94] + error_vector13[95] + error_vector13[96] + error_vector13[97] + error_vector13[98] + error_vector13[99] + error_vector13[100] + error_vector13[101] + error_vector13[102] + error_vector13[103] + error_vector13[104] + error_vector13[105] + error_vector13[106] + error_vector13[107] + error_vector13[108] + error_vector13[109] + error_vector13[110] + error_vector13[111] + error_vector13[112] + error_vector13[113] + error_vector13[114] + error_vector13[115] + error_vector13[116] + error_vector13[117] + error_vector13[118] + error_vector13[119] + error_vector13[120] + error_vector13[121] + error_vector13[122] + error_vector13[123] + error_vector13[124] + error_vector13[125] + error_vector13[126] + error_vector13[127] + error_vector13[128] + error_vector13[129] + error_vector13[130] + error_vector13[131] + error_vector13[132] + error_vector13[133] + error_vector13[134] + error_vector13[135] + error_vector13[136] + error_vector13[137] + error_vector13[138] + error_vector13[139] + error_vector13[140] + error_vector13[141] + error_vector13[142] + error_vector13[143] + error_vector13[144] + error_vector13[145] + error_vector13[146] + error_vector13[147] + error_vector13[148] + error_vector13[149] + error_vector13[150] + error_vector13[151] + error_vector13[152] + error_vector13[153] + error_vector13[154] + error_vector13[155] + error_vector13[156] + error_vector13[157] + error_vector13[158] + error_vector13[159] + error_vector13[160] + error_vector13[161] + error_vector13[162] + error_vector13[163] + error_vector13[164] + error_vector13[165] + error_vector13[166] + error_vector13[167] + error_vector13[168] + error_vector13[169] + error_vector13[170] + error_vector13[171] + error_vector13[172] + error_vector13[173] + error_vector13[174] + error_vector13[175] + error_vector13[176] + error_vector13[177] + error_vector13[178] + error_vector13[179] + error_vector13[180] + error_vector13[181] + error_vector13[182] + error_vector13[183] + error_vector13[184] + error_vector13[185] + error_vector13[186] + error_vector13[187] + error_vector13[188] + error_vector13[189] + error_vector13[190] + error_vector13[191] + error_vector13[192] + error_vector13[193] + error_vector13[194] + error_vector13[195] + error_vector13[196] + error_vector13[197] + error_vector13[198] + error_vector13[199] + error_vector13[200] + error_vector13[201] + error_vector13[202] + error_vector13[203] + error_vector13[204] + error_vector13[205] + error_vector13[206] + error_vector13[207] + error_vector13[208] + error_vector13[209] + error_vector13[210] + error_vector13[211] + error_vector13[212] + error_vector13[213] + error_vector13[214] + error_vector13[215] + error_vector13[216] + error_vector13[217] + error_vector13[218] + error_vector13[219] + error_vector13[220] + error_vector13[221] + error_vector13[222] + error_vector13[223] + error_vector13[224] + error_vector13[225] + error_vector13[226] + error_vector13[227] + error_vector13[228] + error_vector13[229] + error_vector13[230] + error_vector13[231] + error_vector13[232] + error_vector13[233] + error_vector13[234] + error_vector13[235] + error_vector13[236] + error_vector13[237] + error_vector13[238]; 
            errs14 <= error_vector14[0] + error_vector14[1] + error_vector14[2] + error_vector14[3] + error_vector14[4] + error_vector14[5] + error_vector14[6] + error_vector14[7] + error_vector14[8] + error_vector14[9] + error_vector14[10] + error_vector14[11] + error_vector14[12] + error_vector14[13] + error_vector14[14] + error_vector14[15] + error_vector14[16] + error_vector14[17] + error_vector14[18] + error_vector14[19] + error_vector14[20] + error_vector14[21] + error_vector14[22] + error_vector14[23] + error_vector14[24] + error_vector14[25] + error_vector14[26] + error_vector14[27] + error_vector14[28] + error_vector14[29] + error_vector14[30] + error_vector14[31] + error_vector14[32] + error_vector14[33] + error_vector14[34] + error_vector14[35] + error_vector14[36] + error_vector14[37] + error_vector14[38] + error_vector14[39] + error_vector14[40] + error_vector14[41] + error_vector14[42] + error_vector14[43] + error_vector14[44] + error_vector14[45] + error_vector14[46] + error_vector14[47] + error_vector14[48] + error_vector14[49] + error_vector14[50] + error_vector14[51] + error_vector14[52] + error_vector14[53] + error_vector14[54] + error_vector14[55] + error_vector14[56] + error_vector14[57] + error_vector14[58] + error_vector14[59] + error_vector14[60] + error_vector14[61] + error_vector14[62] + error_vector14[63] + error_vector14[64] + error_vector14[65] + error_vector14[66] + error_vector14[67] + error_vector14[68] + error_vector14[69] + error_vector14[70] + error_vector14[71] + error_vector14[72] + error_vector14[73] + error_vector14[74] + error_vector14[75] + error_vector14[76] + error_vector14[77] + error_vector14[78] + error_vector14[79] + error_vector14[80] + error_vector14[81] + error_vector14[82] + error_vector14[83] + error_vector14[84] + error_vector14[85] + error_vector14[86] + error_vector14[87] + error_vector14[88] + error_vector14[89] + error_vector14[90] + error_vector14[91] + error_vector14[92] + error_vector14[93] + error_vector14[94] + error_vector14[95] + error_vector14[96] + error_vector14[97] + error_vector14[98] + error_vector14[99] + error_vector14[100] + error_vector14[101] + error_vector14[102] + error_vector14[103] + error_vector14[104] + error_vector14[105] + error_vector14[106] + error_vector14[107] + error_vector14[108] + error_vector14[109] + error_vector14[110] + error_vector14[111] + error_vector14[112] + error_vector14[113] + error_vector14[114] + error_vector14[115] + error_vector14[116] + error_vector14[117] + error_vector14[118] + error_vector14[119] + error_vector14[120] + error_vector14[121] + error_vector14[122] + error_vector14[123] + error_vector14[124] + error_vector14[125] + error_vector14[126] + error_vector14[127] + error_vector14[128] + error_vector14[129] + error_vector14[130] + error_vector14[131] + error_vector14[132] + error_vector14[133] + error_vector14[134] + error_vector14[135] + error_vector14[136] + error_vector14[137] + error_vector14[138] + error_vector14[139] + error_vector14[140] + error_vector14[141] + error_vector14[142] + error_vector14[143] + error_vector14[144] + error_vector14[145] + error_vector14[146] + error_vector14[147] + error_vector14[148] + error_vector14[149] + error_vector14[150] + error_vector14[151] + error_vector14[152] + error_vector14[153] + error_vector14[154] + error_vector14[155] + error_vector14[156] + error_vector14[157] + error_vector14[158] + error_vector14[159] + error_vector14[160] + error_vector14[161] + error_vector14[162] + error_vector14[163] + error_vector14[164] + error_vector14[165] + error_vector14[166] + error_vector14[167] + error_vector14[168] + error_vector14[169] + error_vector14[170] + error_vector14[171] + error_vector14[172] + error_vector14[173] + error_vector14[174] + error_vector14[175] + error_vector14[176] + error_vector14[177] + error_vector14[178] + error_vector14[179] + error_vector14[180] + error_vector14[181] + error_vector14[182] + error_vector14[183] + error_vector14[184] + error_vector14[185] + error_vector14[186] + error_vector14[187] + error_vector14[188] + error_vector14[189] + error_vector14[190] + error_vector14[191] + error_vector14[192] + error_vector14[193] + error_vector14[194] + error_vector14[195] + error_vector14[196] + error_vector14[197] + error_vector14[198] + error_vector14[199] + error_vector14[200] + error_vector14[201] + error_vector14[202] + error_vector14[203] + error_vector14[204] + error_vector14[205] + error_vector14[206] + error_vector14[207] + error_vector14[208] + error_vector14[209] + error_vector14[210] + error_vector14[211] + error_vector14[212] + error_vector14[213] + error_vector14[214] + error_vector14[215] + error_vector14[216] + error_vector14[217] + error_vector14[218] + error_vector14[219] + error_vector14[220] + error_vector14[221] + error_vector14[222] + error_vector14[223] + error_vector14[224] + error_vector14[225] + error_vector14[226] + error_vector14[227] + error_vector14[228] + error_vector14[229] + error_vector14[230] + error_vector14[231] + error_vector14[232] + error_vector14[233] + error_vector14[234] + error_vector14[235] + error_vector14[236] + error_vector14[237] + error_vector14[238]; 
            errs15 <= error_vector15[0] + error_vector15[1] + error_vector15[2] + error_vector15[3] + error_vector15[4] + error_vector15[5] + error_vector15[6] + error_vector15[7] + error_vector15[8] + error_vector15[9] + error_vector15[10] + error_vector15[11] + error_vector15[12] + error_vector15[13] + error_vector15[14] + error_vector15[15] + error_vector15[16] + error_vector15[17] + error_vector15[18] + error_vector15[19] + error_vector15[20] + error_vector15[21] + error_vector15[22] + error_vector15[23] + error_vector15[24] + error_vector15[25] + error_vector15[26] + error_vector15[27] + error_vector15[28] + error_vector15[29] + error_vector15[30] + error_vector15[31] + error_vector15[32] + error_vector15[33] + error_vector15[34] + error_vector15[35] + error_vector15[36] + error_vector15[37] + error_vector15[38] + error_vector15[39] + error_vector15[40] + error_vector15[41] + error_vector15[42] + error_vector15[43] + error_vector15[44] + error_vector15[45] + error_vector15[46] + error_vector15[47] + error_vector15[48] + error_vector15[49] + error_vector15[50] + error_vector15[51] + error_vector15[52] + error_vector15[53] + error_vector15[54] + error_vector15[55] + error_vector15[56] + error_vector15[57] + error_vector15[58] + error_vector15[59] + error_vector15[60] + error_vector15[61] + error_vector15[62] + error_vector15[63] + error_vector15[64] + error_vector15[65] + error_vector15[66] + error_vector15[67] + error_vector15[68] + error_vector15[69] + error_vector15[70] + error_vector15[71] + error_vector15[72] + error_vector15[73] + error_vector15[74] + error_vector15[75] + error_vector15[76] + error_vector15[77] + error_vector15[78] + error_vector15[79] + error_vector15[80] + error_vector15[81] + error_vector15[82] + error_vector15[83] + error_vector15[84] + error_vector15[85] + error_vector15[86] + error_vector15[87] + error_vector15[88] + error_vector15[89] + error_vector15[90] + error_vector15[91] + error_vector15[92] + error_vector15[93] + error_vector15[94] + error_vector15[95] + error_vector15[96] + error_vector15[97] + error_vector15[98] + error_vector15[99] + error_vector15[100] + error_vector15[101] + error_vector15[102] + error_vector15[103] + error_vector15[104] + error_vector15[105] + error_vector15[106] + error_vector15[107] + error_vector15[108] + error_vector15[109] + error_vector15[110] + error_vector15[111] + error_vector15[112] + error_vector15[113] + error_vector15[114] + error_vector15[115] + error_vector15[116] + error_vector15[117] + error_vector15[118] + error_vector15[119] + error_vector15[120] + error_vector15[121] + error_vector15[122] + error_vector15[123] + error_vector15[124] + error_vector15[125] + error_vector15[126] + error_vector15[127] + error_vector15[128] + error_vector15[129] + error_vector15[130] + error_vector15[131] + error_vector15[132] + error_vector15[133] + error_vector15[134] + error_vector15[135] + error_vector15[136] + error_vector15[137] + error_vector15[138] + error_vector15[139] + error_vector15[140] + error_vector15[141] + error_vector15[142] + error_vector15[143] + error_vector15[144] + error_vector15[145] + error_vector15[146] + error_vector15[147] + error_vector15[148] + error_vector15[149] + error_vector15[150] + error_vector15[151] + error_vector15[152] + error_vector15[153] + error_vector15[154] + error_vector15[155] + error_vector15[156] + error_vector15[157] + error_vector15[158] + error_vector15[159] + error_vector15[160] + error_vector15[161] + error_vector15[162] + error_vector15[163] + error_vector15[164] + error_vector15[165] + error_vector15[166] + error_vector15[167] + error_vector15[168] + error_vector15[169] + error_vector15[170] + error_vector15[171] + error_vector15[172] + error_vector15[173] + error_vector15[174] + error_vector15[175] + error_vector15[176] + error_vector15[177] + error_vector15[178] + error_vector15[179] + error_vector15[180] + error_vector15[181] + error_vector15[182] + error_vector15[183] + error_vector15[184] + error_vector15[185] + error_vector15[186] + error_vector15[187] + error_vector15[188] + error_vector15[189] + error_vector15[190] + error_vector15[191] + error_vector15[192] + error_vector15[193] + error_vector15[194] + error_vector15[195] + error_vector15[196] + error_vector15[197] + error_vector15[198] + error_vector15[199] + error_vector15[200] + error_vector15[201] + error_vector15[202] + error_vector15[203] + error_vector15[204] + error_vector15[205] + error_vector15[206] + error_vector15[207] + error_vector15[208] + error_vector15[209] + error_vector15[210] + error_vector15[211] + error_vector15[212] + error_vector15[213] + error_vector15[214] + error_vector15[215] + error_vector15[216] + error_vector15[217] + error_vector15[218] + error_vector15[219] + error_vector15[220] + error_vector15[221] + error_vector15[222] + error_vector15[223] + error_vector15[224] + error_vector15[225] + error_vector15[226] + error_vector15[227] + error_vector15[228] + error_vector15[229] + error_vector15[230] + error_vector15[231] + error_vector15[232] + error_vector15[233] + error_vector15[234] + error_vector15[235] + error_vector15[236] + error_vector15[237] + error_vector15[238]; 
            errs16 <= error_vector16[0] + error_vector16[1] + error_vector16[2] + error_vector16[3] + error_vector16[4] + error_vector16[5] + error_vector16[6] + error_vector16[7] + error_vector16[8] + error_vector16[9] + error_vector16[10] + error_vector16[11] + error_vector16[12] + error_vector16[13] + error_vector16[14] + error_vector16[15] + error_vector16[16] + error_vector16[17] + error_vector16[18] + error_vector16[19] + error_vector16[20] + error_vector16[21] + error_vector16[22] + error_vector16[23] + error_vector16[24] + error_vector16[25] + error_vector16[26] + error_vector16[27] + error_vector16[28] + error_vector16[29] + error_vector16[30] + error_vector16[31] + error_vector16[32] + error_vector16[33] + error_vector16[34] + error_vector16[35] + error_vector16[36] + error_vector16[37] + error_vector16[38] + error_vector16[39] + error_vector16[40] + error_vector16[41] + error_vector16[42] + error_vector16[43] + error_vector16[44] + error_vector16[45] + error_vector16[46] + error_vector16[47] + error_vector16[48] + error_vector16[49] + error_vector16[50] + error_vector16[51] + error_vector16[52] + error_vector16[53] + error_vector16[54] + error_vector16[55] + error_vector16[56] + error_vector16[57] + error_vector16[58] + error_vector16[59] + error_vector16[60] + error_vector16[61] + error_vector16[62] + error_vector16[63] + error_vector16[64] + error_vector16[65] + error_vector16[66] + error_vector16[67] + error_vector16[68] + error_vector16[69] + error_vector16[70] + error_vector16[71] + error_vector16[72] + error_vector16[73] + error_vector16[74] + error_vector16[75] + error_vector16[76] + error_vector16[77] + error_vector16[78] + error_vector16[79] + error_vector16[80] + error_vector16[81] + error_vector16[82] + error_vector16[83] + error_vector16[84] + error_vector16[85] + error_vector16[86] + error_vector16[87] + error_vector16[88] + error_vector16[89] + error_vector16[90] + error_vector16[91] + error_vector16[92] + error_vector16[93] + error_vector16[94] + error_vector16[95] + error_vector16[96] + error_vector16[97] + error_vector16[98] + error_vector16[99] + error_vector16[100] + error_vector16[101] + error_vector16[102] + error_vector16[103] + error_vector16[104] + error_vector16[105] + error_vector16[106] + error_vector16[107] + error_vector16[108] + error_vector16[109] + error_vector16[110] + error_vector16[111] + error_vector16[112] + error_vector16[113] + error_vector16[114] + error_vector16[115] + error_vector16[116] + error_vector16[117] + error_vector16[118] + error_vector16[119] + error_vector16[120] + error_vector16[121] + error_vector16[122] + error_vector16[123] + error_vector16[124] + error_vector16[125] + error_vector16[126] + error_vector16[127] + error_vector16[128] + error_vector16[129] + error_vector16[130] + error_vector16[131] + error_vector16[132] + error_vector16[133] + error_vector16[134] + error_vector16[135] + error_vector16[136] + error_vector16[137] + error_vector16[138] + error_vector16[139] + error_vector16[140] + error_vector16[141] + error_vector16[142] + error_vector16[143] + error_vector16[144] + error_vector16[145] + error_vector16[146] + error_vector16[147] + error_vector16[148] + error_vector16[149] + error_vector16[150] + error_vector16[151] + error_vector16[152] + error_vector16[153] + error_vector16[154] + error_vector16[155] + error_vector16[156] + error_vector16[157] + error_vector16[158] + error_vector16[159] + error_vector16[160] + error_vector16[161] + error_vector16[162] + error_vector16[163] + error_vector16[164] + error_vector16[165] + error_vector16[166] + error_vector16[167] + error_vector16[168] + error_vector16[169] + error_vector16[170] + error_vector16[171] + error_vector16[172] + error_vector16[173] + error_vector16[174] + error_vector16[175] + error_vector16[176] + error_vector16[177] + error_vector16[178] + error_vector16[179] + error_vector16[180] + error_vector16[181] + error_vector16[182] + error_vector16[183] + error_vector16[184] + error_vector16[185] + error_vector16[186] + error_vector16[187] + error_vector16[188] + error_vector16[189] + error_vector16[190] + error_vector16[191] + error_vector16[192] + error_vector16[193] + error_vector16[194] + error_vector16[195] + error_vector16[196] + error_vector16[197] + error_vector16[198] + error_vector16[199] + error_vector16[200] + error_vector16[201] + error_vector16[202] + error_vector16[203] + error_vector16[204] + error_vector16[205] + error_vector16[206] + error_vector16[207] + error_vector16[208] + error_vector16[209] + error_vector16[210] + error_vector16[211] + error_vector16[212] + error_vector16[213] + error_vector16[214] + error_vector16[215] + error_vector16[216] + error_vector16[217] + error_vector16[218] + error_vector16[219] + error_vector16[220] + error_vector16[221] + error_vector16[222] + error_vector16[223] + error_vector16[224] + error_vector16[225] + error_vector16[226] + error_vector16[227] + error_vector16[228] + error_vector16[229] + error_vector16[230] + error_vector16[231] + error_vector16[232] + error_vector16[233] + error_vector16[234] + error_vector16[235] + error_vector16[236] + error_vector16[237] + error_vector16[238]; 

            if (x == 5'd0) begin
                errs <= errs + errs1 + errs2 + errs3 + errs4 + errs5 + errs6 + errs7 + errs8 + errs9 + errs10 + errs11 + errs12 + errs13 + errs14 + errs15;
            end else
                errs <= errs + errs1 + errs2 + errs3 + errs4 + errs5 + errs6 + errs7 + errs8 + errs9 + errs10 + errs11 + errs12 + errs13 + errs14 + errs15 + errs16;
            
            if ((uncoded_last_iter == 4'd0)&&(uncoded == 1'b0))
                errs_u <= errs_u + errs1_u + errs2_u + errs3_u + errs4_u + errs5_u + errs6_u + errs7_u + errs8_u + errs9_u + errs10_u + errs11_u + errs12_u + errs13_u + errs14_u + errs15_u;
            else
                errs_u <= errs_u + errs1_u + errs2_u + errs3_u + errs4_u + errs5_u + errs6_u + errs7_u + errs8_u + errs9_u + errs10_u + errs11_u + errs12_u + errs13_u + errs14_u + errs15_u + errs16_u;

            if (x == 5'd14)
                sims <= sims + 1;

//            error_vector_u1 <= FIFO_1[(n-1):0] ^ received1;
//            error_vector_u2 <= FIFO_2[(n-1):0] ^ received2;
//            error_vector_u3 <= FIFO_3[(n-1):0] ^ received3;
//            error_vector_u4 <= FIFO_4[(n-1):0] ^ received4;
//            error_vector_u5 <= FIFO_5[(n-1):0] ^ received5;
//            error_vector_u6 <= FIFO_6[(n-1):0] ^ received6;
//            error_vector_u7 <= FIFO_7[(n-1):0] ^ received7;
//            error_vector_u8 <= FIFO_8[(n-1):0] ^ received8;
//            error_vector_u9 <= FIFO_9[(n-1):0] ^ received9;
//            error_vector_u10 <= FIFO_10[(n-1):0] ^ received10;
//            error_vector_u11 <= FIFO_11[(n-1):0] ^ received11;
//            error_vector_u12 <= FIFO_12[(n-1):0] ^ received12;
//            error_vector_u13 <= FIFO_13[(n-1):0] ^ received13;
//            error_vector_u14 <= FIFO_14[(n-1):0] ^ received14;
//            error_vector_u15 <= FIFO_15[(n-1):0] ^ received15;
//            error_vector_u16 <= FIFO_16[(n-1):0] ^ received16;

        end else begin
//            errs_u <= 64'd0;
            fifo_depth <= iterations*16;
            errs <= 64'd0;
            errs_u <= 64'd0;
            counting <= 1'b0;
            sims <= 64'd0;
            valid_err_count <= 1'b0;
            x <= 5'b0;
            uncoded_last_iter <= 4'b0;
            
            error_vector1 <= 0;
            error_vector2 <= 0;
            error_vector3 <= 0;
            error_vector4 <= 0;
            error_vector5 <= 0;
            error_vector6 <= 0;
            error_vector7 <= 0;
            error_vector8 <= 0;
            error_vector9 <= 0;
            error_vector10 <= 0;
            error_vector11 <= 0;
            error_vector12 <= 0;
            error_vector13 <= 0;
            error_vector14 <= 0;
            error_vector15 <= 0;
            error_vector16 <= 0;

            error_u_vector1 <= 0;
            error_u_vector2 <= 0;
            error_u_vector3 <= 0;
            error_u_vector4 <= 0;
            error_u_vector5 <= 0;
            error_u_vector6 <= 0;
            error_u_vector7 <= 0;
            error_u_vector8 <= 0;
            error_u_vector9 <= 0;
            error_u_vector10 <= 0;
            error_u_vector11 <= 0;
            error_u_vector12 <= 0;
            error_u_vector13 <= 0;
            error_u_vector14 <= 0;
            error_u_vector15 <= 0;
            error_u_vector16 <= 0;
            
            errs1 <= 0;
            errs2 <= 0;
            errs3 <= 0;
            errs4 <= 0;
            errs5 <= 0;
            errs6 <= 0;
            errs7 <= 0;
            errs8 <= 0;
            errs9 <= 0;
            errs10 <= 0;
            errs11 <= 0;
            errs12 <= 0;
            errs13 <= 0;
            errs14 <= 0;
            errs15 <= 0;
            errs16 <= 0;

            errs1_u <= 0;
            errs2_u <= 0;
            errs3_u <= 0;
            errs4_u <= 0;
            errs5_u <= 0;
            errs6_u <= 0;
            errs7_u <= 0;
            errs8_u <= 0;
            errs9_u <= 0;
            errs10_u <= 0;
            errs11_u <= 0;
            errs12_u <= 0;
            errs13_u <= 0;
            errs14_u <= 0;
            errs15_u <= 0;
            errs16_u <= 0;
        end
    end
endmodule

