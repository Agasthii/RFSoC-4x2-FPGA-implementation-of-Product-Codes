`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/07/2024 09:06:11 AM
// Design Name: 
// Module Name: PC_decoding_block_ebch_256_239
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PC_decoding_block_ebch_256_239 #(
    parameter n = 256,
    parameter depth = 16
    )(
    input clk,
    input reset,
    input new,
    input [4:0] iter,
    input wire [n-1:0] rec1,
    input wire [n-1:0] rec2,
    input wire [n-1:0] rec3,
    input wire [n-1:0] rec4,
    input wire [n-1:0] rec5,
    input wire [n-1:0] rec6,
    input wire [n-1:0] rec7,
    input wire [n-1:0] rec8,
    input wire [n-1:0] rec9,
    input wire [n-1:0] rec10,
    input wire [n-1:0] rec11,
    input wire [n-1:0] rec12,
    input wire [n-1:0] rec13,
    input wire [n-1:0] rec14,
    input wire [n-1:0] rec15,
    input wire [n-1:0] rec16,
    output reg valid1,
    output reg valid2,
    output reg valid_err,
    output reg hold_enc,
    output reg [n-1:0] dec1,
    output reg [n-1:0] dec2,
    output reg [n-1:0] dec3,
    output reg [n-1:0] dec4,
    output reg [n-1:0] dec5,
    output reg [n-1:0] dec6,
    output reg [n-1:0] dec7,
    output reg [n-1:0] dec8,
    output reg [n-1:0] dec9,
    output reg [n-1:0] dec10,
    output reg [n-1:0] dec11,
    output reg [n-1:0] dec12,
    output reg [n-1:0] dec13,
    output reg [n-1:0] dec14,
    output reg [n-1:0] dec15,
    output reg [n-1:0] dec16
    );
    
    // The control variables
    reg [5:0] counter = 6'b0; 
    reg hold;
    reg [5:0] rounds;
    reg [3:0] C;
    reg temp;
    
    // The inputs to the decoders
    reg [n-1:0] in_rec1;
    reg [n-1:0] in_rec2;
    reg [n-1:0] in_rec3;
    reg [n-1:0] in_rec4;
    reg [n-1:0] in_rec5;
    reg [n-1:0] in_rec6;
    reg [n-1:0] in_rec7;
    reg [n-1:0] in_rec8;
    reg [n-1:0] in_rec9;
    reg [n-1:0] in_rec10;
    reg [n-1:0] in_rec11;
    reg [n-1:0] in_rec12;
    reg [n-1:0] in_rec13;
    reg [n-1:0] in_rec14;
    reg [n-1:0] in_rec15;
    reg [n-1:0] in_rec16;
    
    // The outputs from the decoders
    wire [n-1:0] out_dec1;
    wire [n-1:0] out_dec2;
    wire [n-1:0] out_dec3;
    wire [n-1:0] out_dec4;
    wire [n-1:0] out_dec5;
    wire [n-1:0] out_dec6;
    wire [n-1:0] out_dec7;
    wire [n-1:0] out_dec8;
    wire [n-1:0] out_dec9;
    wire [n-1:0] out_dec10;
    wire [n-1:0] out_dec11;
    wire [n-1:0] out_dec12;
    wire [n-1:0] out_dec13;
    wire [n-1:0] out_dec14;
    wire [n-1:0] out_dec15;
    wire [n-1:0] out_dec16;
    
    // The buffer for the row decoded outputs
    reg [n*depth-1:0] codeword_buf1;
    reg [n*depth-1:0] codeword_buf2;
    reg [n*depth-1:0] codeword_buf3;
    reg [n*depth-1:0] codeword_buf4;
    reg [n*depth-1:0] codeword_buf5;
    reg [n*depth-1:0] codeword_buf6;
    reg [n*depth-1:0] codeword_buf7;
    reg [n*depth-1:0] codeword_buf8;
    reg [n*depth-1:0] codeword_buf9;
    reg [n*depth-1:0] codeword_buf10;
    reg [n*depth-1:0] codeword_buf11;
    reg [n*depth-1:0] codeword_buf12;
    reg [n*depth-1:0] codeword_buf13;
    reg [n*depth-1:0] codeword_buf14;
    reg [n*depth-1:0] codeword_buf15;
    reg [n*depth-1:0] codeword_buf16; 
    
    // The buffer for the col decoded outputs
    reg [n*depth-1:0] codeword_buf2_1;
    reg [n*depth-1:0] codeword_buf2_2;
    reg [n*depth-1:0] codeword_buf2_3;
    reg [n*depth-1:0] codeword_buf2_4;
    reg [n*depth-1:0] codeword_buf2_5;
    reg [n*depth-1:0] codeword_buf2_6;
    reg [n*depth-1:0] codeword_buf2_7;
    reg [n*depth-1:0] codeword_buf2_8;
    reg [n*depth-1:0] codeword_buf2_9;
    reg [n*depth-1:0] codeword_buf2_10;
    reg [n*depth-1:0] codeword_buf2_11;
    reg [n*depth-1:0] codeword_buf2_12;
    reg [n*depth-1:0] codeword_buf2_13;
    reg [n*depth-1:0] codeword_buf2_14;
    reg [n*depth-1:0] codeword_buf2_15;
    reg [n*depth-1:0] codeword_buf2_16; 
    
    bchdecoder_256_239 decoder1(
        .clk(clk),
        .reset(reset),
        .r(in_rec1),
        .dec(out_dec1)
        );
    bchdecoder_256_239 decoder2(
        .clk(clk),
        .reset(reset),
        .r(in_rec2),
        .dec(out_dec2)
        );
    bchdecoder_256_239 decoder3(
        .clk(clk),
        .reset(reset),
        .r(in_rec3),
        .dec(out_dec3)
        );
    bchdecoder_256_239 decoder4(
        .clk(clk),
        .reset(reset),
        .r(in_rec4),
        .dec(out_dec4)
        );
    bchdecoder_256_239 decoder5(
        .clk(clk),
        .reset(reset),
        .r(in_rec5),
        .dec(out_dec5)
        );
    bchdecoder_256_239 decoder6(
        .clk(clk),
        .reset(reset),
        .r(in_rec6),
        .dec(out_dec6)
        );
    bchdecoder_256_239 decoder7(
        .clk(clk),
        .reset(reset),
        .r(in_rec7),
        .dec(out_dec7)
        );
    bchdecoder_256_239 decoder8(
        .clk(clk),
        .reset(reset),
        .r(in_rec8),
        .dec(out_dec8)
        );
    bchdecoder_256_239 decoder9(
        .clk(clk),
        .reset(reset),
        .r(in_rec9),
        .dec(out_dec9)
        );
    bchdecoder_256_239 decoder10(
        .clk(clk),
        .reset(reset),
        .r(in_rec10),
        .dec(out_dec10)
        );
    bchdecoder_256_239 decoder11(
        .clk(clk),
        .reset(reset),
        .r(in_rec11),
        .dec(out_dec11)
        );
    bchdecoder_256_239 decoder12(
        .clk(clk),
        .reset(reset),
        .r(in_rec12),
        .dec(out_dec12)
        );
    bchdecoder_256_239 decoder13(
        .clk(clk),
        .reset(reset),
        .r(in_rec13),
        .dec(out_dec13)
        );
    bchdecoder_256_239 decoder14(
        .clk(clk),
        .reset(reset),
        .r(in_rec14),
        .dec(out_dec14)
        );
    bchdecoder_256_239 decoder15(
        .clk(clk),
        .reset(reset),
        .r(in_rec15),
        .dec(out_dec15)
        );
    bchdecoder_256_239 decoder16(
        .clk(clk),
        .reset(reset),
        .r(in_rec16),
        .dec(out_dec16)
        );
      
    always @(posedge clk) begin
    
        // If the system is ON
        if (reset) begin
            if (new) begin // If New is True
                hold <= 1'b1;
            end
            
            // If the counter value is more than or equal to 41, send the signal to start encoding
            if ((counter >= 6'd29)||(counter <= 6'd12))
                hold_enc <= 1'b1;
            else
                hold_enc <= 1'b0;
                    
            //// Start of the decoding ////
            if (hold) begin // 
            
                //// Start of the row decoding block ////
                if (counter < 6'd23) begin
                
//                    // Encode new codewords if counter vlues is lower than 11
//                    if (counter < 6'd11)    
//                        hold_enc <= 1'b1;
//                    else                
//                        hold_enc <= 1'b0;
                
                    // Give the channel outputs to the row decoder
                    in_rec1  <= rec1;
                    in_rec2  <= rec2;
                    in_rec3  <= rec3;
                    in_rec4  <= rec4;
                    in_rec5  <= rec5;
                    in_rec6  <= rec6;
                    in_rec7  <= rec7;
                    in_rec8  <= rec8;
                    in_rec9  <= rec9;
                    in_rec10 <= rec10;
                    in_rec11 <= rec11;
                    in_rec12 <= rec12;
                    in_rec13 <= rec13;
                    in_rec14 <= rec14;
                    in_rec15 <= rec15;
                    in_rec16 <= rec16;
                    
                    // Shift the row decoded buffer to add the new row decoded outputs
                    codeword_buf1  <= (codeword_buf1  << n);
                    codeword_buf2  <= (codeword_buf2  << n);
                    codeword_buf3  <= (codeword_buf3  << n);
                    codeword_buf4  <= (codeword_buf4  << n);
                    codeword_buf5  <= (codeword_buf5  << n);
                    codeword_buf6  <= (codeword_buf6  << n);
                    codeword_buf7  <= (codeword_buf7  << n);
                    codeword_buf8  <= (codeword_buf8  << n);
                    codeword_buf9  <= (codeword_buf9  << n);
                    codeword_buf10 <= (codeword_buf10 << n);
                    codeword_buf11 <= (codeword_buf11 << n);
                    codeword_buf12 <= (codeword_buf12 << n);
                    codeword_buf13 <= (codeword_buf13 << n);
                    codeword_buf14 <= (codeword_buf14 << n);
                    codeword_buf15 <= (codeword_buf15 << n);
                    codeword_buf16 <= (codeword_buf16 << n);
                    
                    // Put the row decoded outputs to a buffer to be used in col decoding
                    codeword_buf1[(n-1):0]  <= out_dec1;
                    codeword_buf2[(n-1):0]  <= out_dec2;
                    codeword_buf3[(n-1):0]  <= out_dec3;
                    codeword_buf4[(n-1):0]  <= out_dec4;
                    codeword_buf5[(n-1):0]  <= out_dec5;
                    codeword_buf6[(n-1):0]  <= out_dec6;
                    codeword_buf7[(n-1):0]  <= out_dec7;
                    codeword_buf8[(n-1):0]  <= out_dec8;
                    codeword_buf9[(n-1):0]  <= out_dec9;
                    codeword_buf10[(n-1):0] <= out_dec10;
                    codeword_buf11[(n-1):0] <= out_dec11;
                    codeword_buf12[(n-1):0] <= out_dec12;
                    codeword_buf13[(n-1):0] <= out_dec13;
                    codeword_buf14[(n-1):0] <= out_dec14;
                    codeword_buf15[(n-1):0] <= out_dec15;
                    codeword_buf16[(n-1):0] <= out_dec16;
                    
                    // Output x as output because the fully decoded outputs are not yet processed
                    dec1  <= 256'bx;
                    dec2  <= 256'bx;
                    dec3  <= 256'bx;
                    dec4  <= 256'bx;
                    dec5  <= 256'bx;
                    dec6  <= 256'bx;
                    dec7  <= 256'bx;
                    dec8  <= 256'bx;
                    dec9  <= 256'bx;
                    dec10 <= 256'bx;
                    dec11 <= 256'bx;
                    dec12 <= 256'bx;
                    dec13 <= 256'bx;
                    dec14 <= 256'bx;
                    dec15 <= 256'bx;
                    dec16 <= 256'bx;
                    
//                    // Change the valid1
//                    if (counter < 6'd0)
//                        valid1 <= 1'b1;
//                    else
//                        valid1 <= 1'b0;
                    
                    // Increment the counter
                    counter <= counter + 6'b1;
                    
                    // Assign valid2 and valid_err
                    valid2 <= 1'b0;
                    
//                    if ((counter == 6'd0)&&(valid2))
//                        valid_err <= 1'b1;
//                    else
//                        valid_err <= 1'b0;
                    
                    // If the row encoding is done, reduce he rounds count by one, and change C value to 15
                    if (counter == 6'd22) begin 
                        rounds <= rounds - 1;
                        C <= 4'd0;
                    end
                //// End of the row decoding block ////
                
                
                //// Start of the column decoding block //// 
                end else begin
                
                    if (counter < 6'd46) begin
                        // If counter < 39, give the column decoder inputs from the buffer
                        if (counter < 6'd40) begin
                            in_rec1 <= {codeword_buf16[n*0+(16*C+0)],codeword_buf15[n*0+(16*C+0)],codeword_buf14[n*0+(16*C+0)],codeword_buf13[n*0+(16*C+0)],codeword_buf12[n*0+(16*C+0)],codeword_buf11[n*0+(16*C+0)],codeword_buf10[n*0+(16*C+0)],codeword_buf9[n*0+(16*C+0)],codeword_buf8[n*0+(16*C+0)],codeword_buf7[n*0+(16*C+0)],codeword_buf6[n*0+(16*C+0)],codeword_buf5[n*0+(16*C+0)],codeword_buf4[n*0+(16*C+0)],codeword_buf3[n*0+(16*C+0)],codeword_buf2[n*0+(16*C+0)],codeword_buf1[n*0+(16*C+0)],codeword_buf16[n*1+(16*C+0)],codeword_buf15[n*1+(16*C+0)],codeword_buf14[n*1+(16*C+0)],codeword_buf13[n*1+(16*C+0)],codeword_buf12[n*1+(16*C+0)],codeword_buf11[n*1+(16*C+0)],codeword_buf10[n*1+(16*C+0)],codeword_buf9[n*1+(16*C+0)],codeword_buf8[n*1+(16*C+0)],codeword_buf7[n*1+(16*C+0)],codeword_buf6[n*1+(16*C+0)],codeword_buf5[n*1+(16*C+0)],codeword_buf4[n*1+(16*C+0)],codeword_buf3[n*1+(16*C+0)],codeword_buf2[n*1+(16*C+0)],codeword_buf1[n*1+(16*C+0)],codeword_buf16[n*2+(16*C+0)],codeword_buf15[n*2+(16*C+0)],codeword_buf14[n*2+(16*C+0)],codeword_buf13[n*2+(16*C+0)],codeword_buf12[n*2+(16*C+0)],codeword_buf11[n*2+(16*C+0)],codeword_buf10[n*2+(16*C+0)],codeword_buf9[n*2+(16*C+0)],codeword_buf8[n*2+(16*C+0)],codeword_buf7[n*2+(16*C+0)],codeword_buf6[n*2+(16*C+0)],codeword_buf5[n*2+(16*C+0)],codeword_buf4[n*2+(16*C+0)],codeword_buf3[n*2+(16*C+0)],codeword_buf2[n*2+(16*C+0)],codeword_buf1[n*2+(16*C+0)],codeword_buf16[n*3+(16*C+0)],codeword_buf15[n*3+(16*C+0)],codeword_buf14[n*3+(16*C+0)],codeword_buf13[n*3+(16*C+0)],codeword_buf12[n*3+(16*C+0)],codeword_buf11[n*3+(16*C+0)],codeword_buf10[n*3+(16*C+0)],codeword_buf9[n*3+(16*C+0)],codeword_buf8[n*3+(16*C+0)],codeword_buf7[n*3+(16*C+0)],codeword_buf6[n*3+(16*C+0)],codeword_buf5[n*3+(16*C+0)],codeword_buf4[n*3+(16*C+0)],codeword_buf3[n*3+(16*C+0)],codeword_buf2[n*3+(16*C+0)],codeword_buf1[n*3+(16*C+0)],codeword_buf16[n*4+(16*C+0)],codeword_buf15[n*4+(16*C+0)],codeword_buf14[n*4+(16*C+0)],codeword_buf13[n*4+(16*C+0)],codeword_buf12[n*4+(16*C+0)],codeword_buf11[n*4+(16*C+0)],codeword_buf10[n*4+(16*C+0)],codeword_buf9[n*4+(16*C+0)],codeword_buf8[n*4+(16*C+0)],codeword_buf7[n*4+(16*C+0)],codeword_buf6[n*4+(16*C+0)],codeword_buf5[n*4+(16*C+0)],codeword_buf4[n*4+(16*C+0)],codeword_buf3[n*4+(16*C+0)],codeword_buf2[n*4+(16*C+0)],codeword_buf1[n*4+(16*C+0)],codeword_buf16[n*5+(16*C+0)],codeword_buf15[n*5+(16*C+0)],codeword_buf14[n*5+(16*C+0)],codeword_buf13[n*5+(16*C+0)],codeword_buf12[n*5+(16*C+0)],codeword_buf11[n*5+(16*C+0)],codeword_buf10[n*5+(16*C+0)],codeword_buf9[n*5+(16*C+0)],codeword_buf8[n*5+(16*C+0)],codeword_buf7[n*5+(16*C+0)],codeword_buf6[n*5+(16*C+0)],codeword_buf5[n*5+(16*C+0)],codeword_buf4[n*5+(16*C+0)],codeword_buf3[n*5+(16*C+0)],codeword_buf2[n*5+(16*C+0)],codeword_buf1[n*5+(16*C+0)],codeword_buf16[n*6+(16*C+0)],codeword_buf15[n*6+(16*C+0)],codeword_buf14[n*6+(16*C+0)],codeword_buf13[n*6+(16*C+0)],codeword_buf12[n*6+(16*C+0)],codeword_buf11[n*6+(16*C+0)],codeword_buf10[n*6+(16*C+0)],codeword_buf9[n*6+(16*C+0)],codeword_buf8[n*6+(16*C+0)],codeword_buf7[n*6+(16*C+0)],codeword_buf6[n*6+(16*C+0)],codeword_buf5[n*6+(16*C+0)],codeword_buf4[n*6+(16*C+0)],codeword_buf3[n*6+(16*C+0)],codeword_buf2[n*6+(16*C+0)],codeword_buf1[n*6+(16*C+0)],codeword_buf16[n*7+(16*C+0)],codeword_buf15[n*7+(16*C+0)],codeword_buf14[n*7+(16*C+0)],codeword_buf13[n*7+(16*C+0)],codeword_buf12[n*7+(16*C+0)],codeword_buf11[n*7+(16*C+0)],codeword_buf10[n*7+(16*C+0)],codeword_buf9[n*7+(16*C+0)],codeword_buf8[n*7+(16*C+0)],codeword_buf7[n*7+(16*C+0)],codeword_buf6[n*7+(16*C+0)],codeword_buf5[n*7+(16*C+0)],codeword_buf4[n*7+(16*C+0)],codeword_buf3[n*7+(16*C+0)],codeword_buf2[n*7+(16*C+0)],codeword_buf1[n*7+(16*C+0)],codeword_buf16[n*8+(16*C+0)],codeword_buf15[n*8+(16*C+0)],codeword_buf14[n*8+(16*C+0)],codeword_buf13[n*8+(16*C+0)],codeword_buf12[n*8+(16*C+0)],codeword_buf11[n*8+(16*C+0)],codeword_buf10[n*8+(16*C+0)],codeword_buf9[n*8+(16*C+0)],codeword_buf8[n*8+(16*C+0)],codeword_buf7[n*8+(16*C+0)],codeword_buf6[n*8+(16*C+0)],codeword_buf5[n*8+(16*C+0)],codeword_buf4[n*8+(16*C+0)],codeword_buf3[n*8+(16*C+0)],codeword_buf2[n*8+(16*C+0)],codeword_buf1[n*8+(16*C+0)],codeword_buf16[n*9+(16*C+0)],codeword_buf15[n*9+(16*C+0)],codeword_buf14[n*9+(16*C+0)],codeword_buf13[n*9+(16*C+0)],codeword_buf12[n*9+(16*C+0)],codeword_buf11[n*9+(16*C+0)],codeword_buf10[n*9+(16*C+0)],codeword_buf9[n*9+(16*C+0)],codeword_buf8[n*9+(16*C+0)],codeword_buf7[n*9+(16*C+0)],codeword_buf6[n*9+(16*C+0)],codeword_buf5[n*9+(16*C+0)],codeword_buf4[n*9+(16*C+0)],codeword_buf3[n*9+(16*C+0)],codeword_buf2[n*9+(16*C+0)],codeword_buf1[n*9+(16*C+0)],codeword_buf16[n*10+(16*C+0)],codeword_buf15[n*10+(16*C+0)],codeword_buf14[n*10+(16*C+0)],codeword_buf13[n*10+(16*C+0)],codeword_buf12[n*10+(16*C+0)],codeword_buf11[n*10+(16*C+0)],codeword_buf10[n*10+(16*C+0)],codeword_buf9[n*10+(16*C+0)],codeword_buf8[n*10+(16*C+0)],codeword_buf7[n*10+(16*C+0)],codeword_buf6[n*10+(16*C+0)],codeword_buf5[n*10+(16*C+0)],codeword_buf4[n*10+(16*C+0)],codeword_buf3[n*10+(16*C+0)],codeword_buf2[n*10+(16*C+0)],codeword_buf1[n*10+(16*C+0)],codeword_buf16[n*11+(16*C+0)],codeword_buf15[n*11+(16*C+0)],codeword_buf14[n*11+(16*C+0)],codeword_buf13[n*11+(16*C+0)],codeword_buf12[n*11+(16*C+0)],codeword_buf11[n*11+(16*C+0)],codeword_buf10[n*11+(16*C+0)],codeword_buf9[n*11+(16*C+0)],codeword_buf8[n*11+(16*C+0)],codeword_buf7[n*11+(16*C+0)],codeword_buf6[n*11+(16*C+0)],codeword_buf5[n*11+(16*C+0)],codeword_buf4[n*11+(16*C+0)],codeword_buf3[n*11+(16*C+0)],codeword_buf2[n*11+(16*C+0)],codeword_buf1[n*11+(16*C+0)],codeword_buf16[n*12+(16*C+0)],codeword_buf15[n*12+(16*C+0)],codeword_buf14[n*12+(16*C+0)],codeword_buf13[n*12+(16*C+0)],codeword_buf12[n*12+(16*C+0)],codeword_buf11[n*12+(16*C+0)],codeword_buf10[n*12+(16*C+0)],codeword_buf9[n*12+(16*C+0)],codeword_buf8[n*12+(16*C+0)],codeword_buf7[n*12+(16*C+0)],codeword_buf6[n*12+(16*C+0)],codeword_buf5[n*12+(16*C+0)],codeword_buf4[n*12+(16*C+0)],codeword_buf3[n*12+(16*C+0)],codeword_buf2[n*12+(16*C+0)],codeword_buf1[n*12+(16*C+0)],codeword_buf16[n*13+(16*C+0)],codeword_buf15[n*13+(16*C+0)],codeword_buf14[n*13+(16*C+0)],codeword_buf13[n*13+(16*C+0)],codeword_buf12[n*13+(16*C+0)],codeword_buf11[n*13+(16*C+0)],codeword_buf10[n*13+(16*C+0)],codeword_buf9[n*13+(16*C+0)],codeword_buf8[n*13+(16*C+0)],codeword_buf7[n*13+(16*C+0)],codeword_buf6[n*13+(16*C+0)],codeword_buf5[n*13+(16*C+0)],codeword_buf4[n*13+(16*C+0)],codeword_buf3[n*13+(16*C+0)],codeword_buf2[n*13+(16*C+0)],codeword_buf1[n*13+(16*C+0)],codeword_buf16[n*14+(16*C+0)],codeword_buf15[n*14+(16*C+0)],codeword_buf14[n*14+(16*C+0)],codeword_buf13[n*14+(16*C+0)],codeword_buf12[n*14+(16*C+0)],codeword_buf11[n*14+(16*C+0)],codeword_buf10[n*14+(16*C+0)],codeword_buf9[n*14+(16*C+0)],codeword_buf8[n*14+(16*C+0)],codeword_buf7[n*14+(16*C+0)],codeword_buf6[n*14+(16*C+0)],codeword_buf5[n*14+(16*C+0)],codeword_buf4[n*14+(16*C+0)],codeword_buf3[n*14+(16*C+0)],codeword_buf2[n*14+(16*C+0)],codeword_buf1[n*14+(16*C+0)],codeword_buf16[n*15+(16*C+0)],codeword_buf15[n*15+(16*C+0)],codeword_buf14[n*15+(16*C+0)],codeword_buf13[n*15+(16*C+0)],codeword_buf12[n*15+(16*C+0)],codeword_buf11[n*15+(16*C+0)],codeword_buf10[n*15+(16*C+0)],codeword_buf9[n*15+(16*C+0)],codeword_buf8[n*15+(16*C+0)],codeword_buf7[n*15+(16*C+0)],codeword_buf6[n*15+(16*C+0)],codeword_buf5[n*15+(16*C+0)],codeword_buf4[n*15+(16*C+0)],codeword_buf3[n*15+(16*C+0)],codeword_buf2[n*15+(16*C+0)],codeword_buf1[n*15+(16*C+0)]};
                            in_rec2 <= {codeword_buf16[n*0+(16*C+1)],codeword_buf15[n*0+(16*C+1)],codeword_buf14[n*0+(16*C+1)],codeword_buf13[n*0+(16*C+1)],codeword_buf12[n*0+(16*C+1)],codeword_buf11[n*0+(16*C+1)],codeword_buf10[n*0+(16*C+1)],codeword_buf9[n*0+(16*C+1)],codeword_buf8[n*0+(16*C+1)],codeword_buf7[n*0+(16*C+1)],codeword_buf6[n*0+(16*C+1)],codeword_buf5[n*0+(16*C+1)],codeword_buf4[n*0+(16*C+1)],codeword_buf3[n*0+(16*C+1)],codeword_buf2[n*0+(16*C+1)],codeword_buf1[n*0+(16*C+1)],codeword_buf16[n*1+(16*C+1)],codeword_buf15[n*1+(16*C+1)],codeword_buf14[n*1+(16*C+1)],codeword_buf13[n*1+(16*C+1)],codeword_buf12[n*1+(16*C+1)],codeword_buf11[n*1+(16*C+1)],codeword_buf10[n*1+(16*C+1)],codeword_buf9[n*1+(16*C+1)],codeword_buf8[n*1+(16*C+1)],codeword_buf7[n*1+(16*C+1)],codeword_buf6[n*1+(16*C+1)],codeword_buf5[n*1+(16*C+1)],codeword_buf4[n*1+(16*C+1)],codeword_buf3[n*1+(16*C+1)],codeword_buf2[n*1+(16*C+1)],codeword_buf1[n*1+(16*C+1)],codeword_buf16[n*2+(16*C+1)],codeword_buf15[n*2+(16*C+1)],codeword_buf14[n*2+(16*C+1)],codeword_buf13[n*2+(16*C+1)],codeword_buf12[n*2+(16*C+1)],codeword_buf11[n*2+(16*C+1)],codeword_buf10[n*2+(16*C+1)],codeword_buf9[n*2+(16*C+1)],codeword_buf8[n*2+(16*C+1)],codeword_buf7[n*2+(16*C+1)],codeword_buf6[n*2+(16*C+1)],codeword_buf5[n*2+(16*C+1)],codeword_buf4[n*2+(16*C+1)],codeword_buf3[n*2+(16*C+1)],codeword_buf2[n*2+(16*C+1)],codeword_buf1[n*2+(16*C+1)],codeword_buf16[n*3+(16*C+1)],codeword_buf15[n*3+(16*C+1)],codeword_buf14[n*3+(16*C+1)],codeword_buf13[n*3+(16*C+1)],codeword_buf12[n*3+(16*C+1)],codeword_buf11[n*3+(16*C+1)],codeword_buf10[n*3+(16*C+1)],codeword_buf9[n*3+(16*C+1)],codeword_buf8[n*3+(16*C+1)],codeword_buf7[n*3+(16*C+1)],codeword_buf6[n*3+(16*C+1)],codeword_buf5[n*3+(16*C+1)],codeword_buf4[n*3+(16*C+1)],codeword_buf3[n*3+(16*C+1)],codeword_buf2[n*3+(16*C+1)],codeword_buf1[n*3+(16*C+1)],codeword_buf16[n*4+(16*C+1)],codeword_buf15[n*4+(16*C+1)],codeword_buf14[n*4+(16*C+1)],codeword_buf13[n*4+(16*C+1)],codeword_buf12[n*4+(16*C+1)],codeword_buf11[n*4+(16*C+1)],codeword_buf10[n*4+(16*C+1)],codeword_buf9[n*4+(16*C+1)],codeword_buf8[n*4+(16*C+1)],codeword_buf7[n*4+(16*C+1)],codeword_buf6[n*4+(16*C+1)],codeword_buf5[n*4+(16*C+1)],codeword_buf4[n*4+(16*C+1)],codeword_buf3[n*4+(16*C+1)],codeword_buf2[n*4+(16*C+1)],codeword_buf1[n*4+(16*C+1)],codeword_buf16[n*5+(16*C+1)],codeword_buf15[n*5+(16*C+1)],codeword_buf14[n*5+(16*C+1)],codeword_buf13[n*5+(16*C+1)],codeword_buf12[n*5+(16*C+1)],codeword_buf11[n*5+(16*C+1)],codeword_buf10[n*5+(16*C+1)],codeword_buf9[n*5+(16*C+1)],codeword_buf8[n*5+(16*C+1)],codeword_buf7[n*5+(16*C+1)],codeword_buf6[n*5+(16*C+1)],codeword_buf5[n*5+(16*C+1)],codeword_buf4[n*5+(16*C+1)],codeword_buf3[n*5+(16*C+1)],codeword_buf2[n*5+(16*C+1)],codeword_buf1[n*5+(16*C+1)],codeword_buf16[n*6+(16*C+1)],codeword_buf15[n*6+(16*C+1)],codeword_buf14[n*6+(16*C+1)],codeword_buf13[n*6+(16*C+1)],codeword_buf12[n*6+(16*C+1)],codeword_buf11[n*6+(16*C+1)],codeword_buf10[n*6+(16*C+1)],codeword_buf9[n*6+(16*C+1)],codeword_buf8[n*6+(16*C+1)],codeword_buf7[n*6+(16*C+1)],codeword_buf6[n*6+(16*C+1)],codeword_buf5[n*6+(16*C+1)],codeword_buf4[n*6+(16*C+1)],codeword_buf3[n*6+(16*C+1)],codeword_buf2[n*6+(16*C+1)],codeword_buf1[n*6+(16*C+1)],codeword_buf16[n*7+(16*C+1)],codeword_buf15[n*7+(16*C+1)],codeword_buf14[n*7+(16*C+1)],codeword_buf13[n*7+(16*C+1)],codeword_buf12[n*7+(16*C+1)],codeword_buf11[n*7+(16*C+1)],codeword_buf10[n*7+(16*C+1)],codeword_buf9[n*7+(16*C+1)],codeword_buf8[n*7+(16*C+1)],codeword_buf7[n*7+(16*C+1)],codeword_buf6[n*7+(16*C+1)],codeword_buf5[n*7+(16*C+1)],codeword_buf4[n*7+(16*C+1)],codeword_buf3[n*7+(16*C+1)],codeword_buf2[n*7+(16*C+1)],codeword_buf1[n*7+(16*C+1)],codeword_buf16[n*8+(16*C+1)],codeword_buf15[n*8+(16*C+1)],codeword_buf14[n*8+(16*C+1)],codeword_buf13[n*8+(16*C+1)],codeword_buf12[n*8+(16*C+1)],codeword_buf11[n*8+(16*C+1)],codeword_buf10[n*8+(16*C+1)],codeword_buf9[n*8+(16*C+1)],codeword_buf8[n*8+(16*C+1)],codeword_buf7[n*8+(16*C+1)],codeword_buf6[n*8+(16*C+1)],codeword_buf5[n*8+(16*C+1)],codeword_buf4[n*8+(16*C+1)],codeword_buf3[n*8+(16*C+1)],codeword_buf2[n*8+(16*C+1)],codeword_buf1[n*8+(16*C+1)],codeword_buf16[n*9+(16*C+1)],codeword_buf15[n*9+(16*C+1)],codeword_buf14[n*9+(16*C+1)],codeword_buf13[n*9+(16*C+1)],codeword_buf12[n*9+(16*C+1)],codeword_buf11[n*9+(16*C+1)],codeword_buf10[n*9+(16*C+1)],codeword_buf9[n*9+(16*C+1)],codeword_buf8[n*9+(16*C+1)],codeword_buf7[n*9+(16*C+1)],codeword_buf6[n*9+(16*C+1)],codeword_buf5[n*9+(16*C+1)],codeword_buf4[n*9+(16*C+1)],codeword_buf3[n*9+(16*C+1)],codeword_buf2[n*9+(16*C+1)],codeword_buf1[n*9+(16*C+1)],codeword_buf16[n*10+(16*C+1)],codeword_buf15[n*10+(16*C+1)],codeword_buf14[n*10+(16*C+1)],codeword_buf13[n*10+(16*C+1)],codeword_buf12[n*10+(16*C+1)],codeword_buf11[n*10+(16*C+1)],codeword_buf10[n*10+(16*C+1)],codeword_buf9[n*10+(16*C+1)],codeword_buf8[n*10+(16*C+1)],codeword_buf7[n*10+(16*C+1)],codeword_buf6[n*10+(16*C+1)],codeword_buf5[n*10+(16*C+1)],codeword_buf4[n*10+(16*C+1)],codeword_buf3[n*10+(16*C+1)],codeword_buf2[n*10+(16*C+1)],codeword_buf1[n*10+(16*C+1)],codeword_buf16[n*11+(16*C+1)],codeword_buf15[n*11+(16*C+1)],codeword_buf14[n*11+(16*C+1)],codeword_buf13[n*11+(16*C+1)],codeword_buf12[n*11+(16*C+1)],codeword_buf11[n*11+(16*C+1)],codeword_buf10[n*11+(16*C+1)],codeword_buf9[n*11+(16*C+1)],codeword_buf8[n*11+(16*C+1)],codeword_buf7[n*11+(16*C+1)],codeword_buf6[n*11+(16*C+1)],codeword_buf5[n*11+(16*C+1)],codeword_buf4[n*11+(16*C+1)],codeword_buf3[n*11+(16*C+1)],codeword_buf2[n*11+(16*C+1)],codeword_buf1[n*11+(16*C+1)],codeword_buf16[n*12+(16*C+1)],codeword_buf15[n*12+(16*C+1)],codeword_buf14[n*12+(16*C+1)],codeword_buf13[n*12+(16*C+1)],codeword_buf12[n*12+(16*C+1)],codeword_buf11[n*12+(16*C+1)],codeword_buf10[n*12+(16*C+1)],codeword_buf9[n*12+(16*C+1)],codeword_buf8[n*12+(16*C+1)],codeword_buf7[n*12+(16*C+1)],codeword_buf6[n*12+(16*C+1)],codeword_buf5[n*12+(16*C+1)],codeword_buf4[n*12+(16*C+1)],codeword_buf3[n*12+(16*C+1)],codeword_buf2[n*12+(16*C+1)],codeword_buf1[n*12+(16*C+1)],codeword_buf16[n*13+(16*C+1)],codeword_buf15[n*13+(16*C+1)],codeword_buf14[n*13+(16*C+1)],codeword_buf13[n*13+(16*C+1)],codeword_buf12[n*13+(16*C+1)],codeword_buf11[n*13+(16*C+1)],codeword_buf10[n*13+(16*C+1)],codeword_buf9[n*13+(16*C+1)],codeword_buf8[n*13+(16*C+1)],codeword_buf7[n*13+(16*C+1)],codeword_buf6[n*13+(16*C+1)],codeword_buf5[n*13+(16*C+1)],codeword_buf4[n*13+(16*C+1)],codeword_buf3[n*13+(16*C+1)],codeword_buf2[n*13+(16*C+1)],codeword_buf1[n*13+(16*C+1)],codeword_buf16[n*14+(16*C+1)],codeword_buf15[n*14+(16*C+1)],codeword_buf14[n*14+(16*C+1)],codeword_buf13[n*14+(16*C+1)],codeword_buf12[n*14+(16*C+1)],codeword_buf11[n*14+(16*C+1)],codeword_buf10[n*14+(16*C+1)],codeword_buf9[n*14+(16*C+1)],codeword_buf8[n*14+(16*C+1)],codeword_buf7[n*14+(16*C+1)],codeword_buf6[n*14+(16*C+1)],codeword_buf5[n*14+(16*C+1)],codeword_buf4[n*14+(16*C+1)],codeword_buf3[n*14+(16*C+1)],codeword_buf2[n*14+(16*C+1)],codeword_buf1[n*14+(16*C+1)],codeword_buf16[n*15+(16*C+1)],codeword_buf15[n*15+(16*C+1)],codeword_buf14[n*15+(16*C+1)],codeword_buf13[n*15+(16*C+1)],codeword_buf12[n*15+(16*C+1)],codeword_buf11[n*15+(16*C+1)],codeword_buf10[n*15+(16*C+1)],codeword_buf9[n*15+(16*C+1)],codeword_buf8[n*15+(16*C+1)],codeword_buf7[n*15+(16*C+1)],codeword_buf6[n*15+(16*C+1)],codeword_buf5[n*15+(16*C+1)],codeword_buf4[n*15+(16*C+1)],codeword_buf3[n*15+(16*C+1)],codeword_buf2[n*15+(16*C+1)],codeword_buf1[n*15+(16*C+1)]};
                            in_rec3 <= {codeword_buf16[n*0+(16*C+2)],codeword_buf15[n*0+(16*C+2)],codeword_buf14[n*0+(16*C+2)],codeword_buf13[n*0+(16*C+2)],codeword_buf12[n*0+(16*C+2)],codeword_buf11[n*0+(16*C+2)],codeword_buf10[n*0+(16*C+2)],codeword_buf9[n*0+(16*C+2)],codeword_buf8[n*0+(16*C+2)],codeword_buf7[n*0+(16*C+2)],codeword_buf6[n*0+(16*C+2)],codeword_buf5[n*0+(16*C+2)],codeword_buf4[n*0+(16*C+2)],codeword_buf3[n*0+(16*C+2)],codeword_buf2[n*0+(16*C+2)],codeword_buf1[n*0+(16*C+2)],codeword_buf16[n*1+(16*C+2)],codeword_buf15[n*1+(16*C+2)],codeword_buf14[n*1+(16*C+2)],codeword_buf13[n*1+(16*C+2)],codeword_buf12[n*1+(16*C+2)],codeword_buf11[n*1+(16*C+2)],codeword_buf10[n*1+(16*C+2)],codeword_buf9[n*1+(16*C+2)],codeword_buf8[n*1+(16*C+2)],codeword_buf7[n*1+(16*C+2)],codeword_buf6[n*1+(16*C+2)],codeword_buf5[n*1+(16*C+2)],codeword_buf4[n*1+(16*C+2)],codeword_buf3[n*1+(16*C+2)],codeword_buf2[n*1+(16*C+2)],codeword_buf1[n*1+(16*C+2)],codeword_buf16[n*2+(16*C+2)],codeword_buf15[n*2+(16*C+2)],codeword_buf14[n*2+(16*C+2)],codeword_buf13[n*2+(16*C+2)],codeword_buf12[n*2+(16*C+2)],codeword_buf11[n*2+(16*C+2)],codeword_buf10[n*2+(16*C+2)],codeword_buf9[n*2+(16*C+2)],codeword_buf8[n*2+(16*C+2)],codeword_buf7[n*2+(16*C+2)],codeword_buf6[n*2+(16*C+2)],codeword_buf5[n*2+(16*C+2)],codeword_buf4[n*2+(16*C+2)],codeword_buf3[n*2+(16*C+2)],codeword_buf2[n*2+(16*C+2)],codeword_buf1[n*2+(16*C+2)],codeword_buf16[n*3+(16*C+2)],codeword_buf15[n*3+(16*C+2)],codeword_buf14[n*3+(16*C+2)],codeword_buf13[n*3+(16*C+2)],codeword_buf12[n*3+(16*C+2)],codeword_buf11[n*3+(16*C+2)],codeword_buf10[n*3+(16*C+2)],codeword_buf9[n*3+(16*C+2)],codeword_buf8[n*3+(16*C+2)],codeword_buf7[n*3+(16*C+2)],codeword_buf6[n*3+(16*C+2)],codeword_buf5[n*3+(16*C+2)],codeword_buf4[n*3+(16*C+2)],codeword_buf3[n*3+(16*C+2)],codeword_buf2[n*3+(16*C+2)],codeword_buf1[n*3+(16*C+2)],codeword_buf16[n*4+(16*C+2)],codeword_buf15[n*4+(16*C+2)],codeword_buf14[n*4+(16*C+2)],codeword_buf13[n*4+(16*C+2)],codeword_buf12[n*4+(16*C+2)],codeword_buf11[n*4+(16*C+2)],codeword_buf10[n*4+(16*C+2)],codeword_buf9[n*4+(16*C+2)],codeword_buf8[n*4+(16*C+2)],codeword_buf7[n*4+(16*C+2)],codeword_buf6[n*4+(16*C+2)],codeword_buf5[n*4+(16*C+2)],codeword_buf4[n*4+(16*C+2)],codeword_buf3[n*4+(16*C+2)],codeword_buf2[n*4+(16*C+2)],codeword_buf1[n*4+(16*C+2)],codeword_buf16[n*5+(16*C+2)],codeword_buf15[n*5+(16*C+2)],codeword_buf14[n*5+(16*C+2)],codeword_buf13[n*5+(16*C+2)],codeword_buf12[n*5+(16*C+2)],codeword_buf11[n*5+(16*C+2)],codeword_buf10[n*5+(16*C+2)],codeword_buf9[n*5+(16*C+2)],codeword_buf8[n*5+(16*C+2)],codeword_buf7[n*5+(16*C+2)],codeword_buf6[n*5+(16*C+2)],codeword_buf5[n*5+(16*C+2)],codeword_buf4[n*5+(16*C+2)],codeword_buf3[n*5+(16*C+2)],codeword_buf2[n*5+(16*C+2)],codeword_buf1[n*5+(16*C+2)],codeword_buf16[n*6+(16*C+2)],codeword_buf15[n*6+(16*C+2)],codeword_buf14[n*6+(16*C+2)],codeword_buf13[n*6+(16*C+2)],codeword_buf12[n*6+(16*C+2)],codeword_buf11[n*6+(16*C+2)],codeword_buf10[n*6+(16*C+2)],codeword_buf9[n*6+(16*C+2)],codeword_buf8[n*6+(16*C+2)],codeword_buf7[n*6+(16*C+2)],codeword_buf6[n*6+(16*C+2)],codeword_buf5[n*6+(16*C+2)],codeword_buf4[n*6+(16*C+2)],codeword_buf3[n*6+(16*C+2)],codeword_buf2[n*6+(16*C+2)],codeword_buf1[n*6+(16*C+2)],codeword_buf16[n*7+(16*C+2)],codeword_buf15[n*7+(16*C+2)],codeword_buf14[n*7+(16*C+2)],codeword_buf13[n*7+(16*C+2)],codeword_buf12[n*7+(16*C+2)],codeword_buf11[n*7+(16*C+2)],codeword_buf10[n*7+(16*C+2)],codeword_buf9[n*7+(16*C+2)],codeword_buf8[n*7+(16*C+2)],codeword_buf7[n*7+(16*C+2)],codeword_buf6[n*7+(16*C+2)],codeword_buf5[n*7+(16*C+2)],codeword_buf4[n*7+(16*C+2)],codeword_buf3[n*7+(16*C+2)],codeword_buf2[n*7+(16*C+2)],codeword_buf1[n*7+(16*C+2)],codeword_buf16[n*8+(16*C+2)],codeword_buf15[n*8+(16*C+2)],codeword_buf14[n*8+(16*C+2)],codeword_buf13[n*8+(16*C+2)],codeword_buf12[n*8+(16*C+2)],codeword_buf11[n*8+(16*C+2)],codeword_buf10[n*8+(16*C+2)],codeword_buf9[n*8+(16*C+2)],codeword_buf8[n*8+(16*C+2)],codeword_buf7[n*8+(16*C+2)],codeword_buf6[n*8+(16*C+2)],codeword_buf5[n*8+(16*C+2)],codeword_buf4[n*8+(16*C+2)],codeword_buf3[n*8+(16*C+2)],codeword_buf2[n*8+(16*C+2)],codeword_buf1[n*8+(16*C+2)],codeword_buf16[n*9+(16*C+2)],codeword_buf15[n*9+(16*C+2)],codeword_buf14[n*9+(16*C+2)],codeword_buf13[n*9+(16*C+2)],codeword_buf12[n*9+(16*C+2)],codeword_buf11[n*9+(16*C+2)],codeword_buf10[n*9+(16*C+2)],codeword_buf9[n*9+(16*C+2)],codeword_buf8[n*9+(16*C+2)],codeword_buf7[n*9+(16*C+2)],codeword_buf6[n*9+(16*C+2)],codeword_buf5[n*9+(16*C+2)],codeword_buf4[n*9+(16*C+2)],codeword_buf3[n*9+(16*C+2)],codeword_buf2[n*9+(16*C+2)],codeword_buf1[n*9+(16*C+2)],codeword_buf16[n*10+(16*C+2)],codeword_buf15[n*10+(16*C+2)],codeword_buf14[n*10+(16*C+2)],codeword_buf13[n*10+(16*C+2)],codeword_buf12[n*10+(16*C+2)],codeword_buf11[n*10+(16*C+2)],codeword_buf10[n*10+(16*C+2)],codeword_buf9[n*10+(16*C+2)],codeword_buf8[n*10+(16*C+2)],codeword_buf7[n*10+(16*C+2)],codeword_buf6[n*10+(16*C+2)],codeword_buf5[n*10+(16*C+2)],codeword_buf4[n*10+(16*C+2)],codeword_buf3[n*10+(16*C+2)],codeword_buf2[n*10+(16*C+2)],codeword_buf1[n*10+(16*C+2)],codeword_buf16[n*11+(16*C+2)],codeword_buf15[n*11+(16*C+2)],codeword_buf14[n*11+(16*C+2)],codeword_buf13[n*11+(16*C+2)],codeword_buf12[n*11+(16*C+2)],codeword_buf11[n*11+(16*C+2)],codeword_buf10[n*11+(16*C+2)],codeword_buf9[n*11+(16*C+2)],codeword_buf8[n*11+(16*C+2)],codeword_buf7[n*11+(16*C+2)],codeword_buf6[n*11+(16*C+2)],codeword_buf5[n*11+(16*C+2)],codeword_buf4[n*11+(16*C+2)],codeword_buf3[n*11+(16*C+2)],codeword_buf2[n*11+(16*C+2)],codeword_buf1[n*11+(16*C+2)],codeword_buf16[n*12+(16*C+2)],codeword_buf15[n*12+(16*C+2)],codeword_buf14[n*12+(16*C+2)],codeword_buf13[n*12+(16*C+2)],codeword_buf12[n*12+(16*C+2)],codeword_buf11[n*12+(16*C+2)],codeword_buf10[n*12+(16*C+2)],codeword_buf9[n*12+(16*C+2)],codeword_buf8[n*12+(16*C+2)],codeword_buf7[n*12+(16*C+2)],codeword_buf6[n*12+(16*C+2)],codeword_buf5[n*12+(16*C+2)],codeword_buf4[n*12+(16*C+2)],codeword_buf3[n*12+(16*C+2)],codeword_buf2[n*12+(16*C+2)],codeword_buf1[n*12+(16*C+2)],codeword_buf16[n*13+(16*C+2)],codeword_buf15[n*13+(16*C+2)],codeword_buf14[n*13+(16*C+2)],codeword_buf13[n*13+(16*C+2)],codeword_buf12[n*13+(16*C+2)],codeword_buf11[n*13+(16*C+2)],codeword_buf10[n*13+(16*C+2)],codeword_buf9[n*13+(16*C+2)],codeword_buf8[n*13+(16*C+2)],codeword_buf7[n*13+(16*C+2)],codeword_buf6[n*13+(16*C+2)],codeword_buf5[n*13+(16*C+2)],codeword_buf4[n*13+(16*C+2)],codeword_buf3[n*13+(16*C+2)],codeword_buf2[n*13+(16*C+2)],codeword_buf1[n*13+(16*C+2)],codeword_buf16[n*14+(16*C+2)],codeword_buf15[n*14+(16*C+2)],codeword_buf14[n*14+(16*C+2)],codeword_buf13[n*14+(16*C+2)],codeword_buf12[n*14+(16*C+2)],codeword_buf11[n*14+(16*C+2)],codeword_buf10[n*14+(16*C+2)],codeword_buf9[n*14+(16*C+2)],codeword_buf8[n*14+(16*C+2)],codeword_buf7[n*14+(16*C+2)],codeword_buf6[n*14+(16*C+2)],codeword_buf5[n*14+(16*C+2)],codeword_buf4[n*14+(16*C+2)],codeword_buf3[n*14+(16*C+2)],codeword_buf2[n*14+(16*C+2)],codeword_buf1[n*14+(16*C+2)],codeword_buf16[n*15+(16*C+2)],codeword_buf15[n*15+(16*C+2)],codeword_buf14[n*15+(16*C+2)],codeword_buf13[n*15+(16*C+2)],codeword_buf12[n*15+(16*C+2)],codeword_buf11[n*15+(16*C+2)],codeword_buf10[n*15+(16*C+2)],codeword_buf9[n*15+(16*C+2)],codeword_buf8[n*15+(16*C+2)],codeword_buf7[n*15+(16*C+2)],codeword_buf6[n*15+(16*C+2)],codeword_buf5[n*15+(16*C+2)],codeword_buf4[n*15+(16*C+2)],codeword_buf3[n*15+(16*C+2)],codeword_buf2[n*15+(16*C+2)],codeword_buf1[n*15+(16*C+2)]};
                            in_rec4 <= {codeword_buf16[n*0+(16*C+3)],codeword_buf15[n*0+(16*C+3)],codeword_buf14[n*0+(16*C+3)],codeword_buf13[n*0+(16*C+3)],codeword_buf12[n*0+(16*C+3)],codeword_buf11[n*0+(16*C+3)],codeword_buf10[n*0+(16*C+3)],codeword_buf9[n*0+(16*C+3)],codeword_buf8[n*0+(16*C+3)],codeword_buf7[n*0+(16*C+3)],codeword_buf6[n*0+(16*C+3)],codeword_buf5[n*0+(16*C+3)],codeword_buf4[n*0+(16*C+3)],codeword_buf3[n*0+(16*C+3)],codeword_buf2[n*0+(16*C+3)],codeword_buf1[n*0+(16*C+3)],codeword_buf16[n*1+(16*C+3)],codeword_buf15[n*1+(16*C+3)],codeword_buf14[n*1+(16*C+3)],codeword_buf13[n*1+(16*C+3)],codeword_buf12[n*1+(16*C+3)],codeword_buf11[n*1+(16*C+3)],codeword_buf10[n*1+(16*C+3)],codeword_buf9[n*1+(16*C+3)],codeword_buf8[n*1+(16*C+3)],codeword_buf7[n*1+(16*C+3)],codeword_buf6[n*1+(16*C+3)],codeword_buf5[n*1+(16*C+3)],codeword_buf4[n*1+(16*C+3)],codeword_buf3[n*1+(16*C+3)],codeword_buf2[n*1+(16*C+3)],codeword_buf1[n*1+(16*C+3)],codeword_buf16[n*2+(16*C+3)],codeword_buf15[n*2+(16*C+3)],codeword_buf14[n*2+(16*C+3)],codeword_buf13[n*2+(16*C+3)],codeword_buf12[n*2+(16*C+3)],codeword_buf11[n*2+(16*C+3)],codeword_buf10[n*2+(16*C+3)],codeword_buf9[n*2+(16*C+3)],codeword_buf8[n*2+(16*C+3)],codeword_buf7[n*2+(16*C+3)],codeword_buf6[n*2+(16*C+3)],codeword_buf5[n*2+(16*C+3)],codeword_buf4[n*2+(16*C+3)],codeword_buf3[n*2+(16*C+3)],codeword_buf2[n*2+(16*C+3)],codeword_buf1[n*2+(16*C+3)],codeword_buf16[n*3+(16*C+3)],codeword_buf15[n*3+(16*C+3)],codeword_buf14[n*3+(16*C+3)],codeword_buf13[n*3+(16*C+3)],codeword_buf12[n*3+(16*C+3)],codeword_buf11[n*3+(16*C+3)],codeword_buf10[n*3+(16*C+3)],codeword_buf9[n*3+(16*C+3)],codeword_buf8[n*3+(16*C+3)],codeword_buf7[n*3+(16*C+3)],codeword_buf6[n*3+(16*C+3)],codeword_buf5[n*3+(16*C+3)],codeword_buf4[n*3+(16*C+3)],codeword_buf3[n*3+(16*C+3)],codeword_buf2[n*3+(16*C+3)],codeword_buf1[n*3+(16*C+3)],codeword_buf16[n*4+(16*C+3)],codeword_buf15[n*4+(16*C+3)],codeword_buf14[n*4+(16*C+3)],codeword_buf13[n*4+(16*C+3)],codeword_buf12[n*4+(16*C+3)],codeword_buf11[n*4+(16*C+3)],codeword_buf10[n*4+(16*C+3)],codeword_buf9[n*4+(16*C+3)],codeword_buf8[n*4+(16*C+3)],codeword_buf7[n*4+(16*C+3)],codeword_buf6[n*4+(16*C+3)],codeword_buf5[n*4+(16*C+3)],codeword_buf4[n*4+(16*C+3)],codeword_buf3[n*4+(16*C+3)],codeword_buf2[n*4+(16*C+3)],codeword_buf1[n*4+(16*C+3)],codeword_buf16[n*5+(16*C+3)],codeword_buf15[n*5+(16*C+3)],codeword_buf14[n*5+(16*C+3)],codeword_buf13[n*5+(16*C+3)],codeword_buf12[n*5+(16*C+3)],codeword_buf11[n*5+(16*C+3)],codeword_buf10[n*5+(16*C+3)],codeword_buf9[n*5+(16*C+3)],codeword_buf8[n*5+(16*C+3)],codeword_buf7[n*5+(16*C+3)],codeword_buf6[n*5+(16*C+3)],codeword_buf5[n*5+(16*C+3)],codeword_buf4[n*5+(16*C+3)],codeword_buf3[n*5+(16*C+3)],codeword_buf2[n*5+(16*C+3)],codeword_buf1[n*5+(16*C+3)],codeword_buf16[n*6+(16*C+3)],codeword_buf15[n*6+(16*C+3)],codeword_buf14[n*6+(16*C+3)],codeword_buf13[n*6+(16*C+3)],codeword_buf12[n*6+(16*C+3)],codeword_buf11[n*6+(16*C+3)],codeword_buf10[n*6+(16*C+3)],codeword_buf9[n*6+(16*C+3)],codeword_buf8[n*6+(16*C+3)],codeword_buf7[n*6+(16*C+3)],codeword_buf6[n*6+(16*C+3)],codeword_buf5[n*6+(16*C+3)],codeword_buf4[n*6+(16*C+3)],codeword_buf3[n*6+(16*C+3)],codeword_buf2[n*6+(16*C+3)],codeword_buf1[n*6+(16*C+3)],codeword_buf16[n*7+(16*C+3)],codeword_buf15[n*7+(16*C+3)],codeword_buf14[n*7+(16*C+3)],codeword_buf13[n*7+(16*C+3)],codeword_buf12[n*7+(16*C+3)],codeword_buf11[n*7+(16*C+3)],codeword_buf10[n*7+(16*C+3)],codeword_buf9[n*7+(16*C+3)],codeword_buf8[n*7+(16*C+3)],codeword_buf7[n*7+(16*C+3)],codeword_buf6[n*7+(16*C+3)],codeword_buf5[n*7+(16*C+3)],codeword_buf4[n*7+(16*C+3)],codeword_buf3[n*7+(16*C+3)],codeword_buf2[n*7+(16*C+3)],codeword_buf1[n*7+(16*C+3)],codeword_buf16[n*8+(16*C+3)],codeword_buf15[n*8+(16*C+3)],codeword_buf14[n*8+(16*C+3)],codeword_buf13[n*8+(16*C+3)],codeword_buf12[n*8+(16*C+3)],codeword_buf11[n*8+(16*C+3)],codeword_buf10[n*8+(16*C+3)],codeword_buf9[n*8+(16*C+3)],codeword_buf8[n*8+(16*C+3)],codeword_buf7[n*8+(16*C+3)],codeword_buf6[n*8+(16*C+3)],codeword_buf5[n*8+(16*C+3)],codeword_buf4[n*8+(16*C+3)],codeword_buf3[n*8+(16*C+3)],codeword_buf2[n*8+(16*C+3)],codeword_buf1[n*8+(16*C+3)],codeword_buf16[n*9+(16*C+3)],codeword_buf15[n*9+(16*C+3)],codeword_buf14[n*9+(16*C+3)],codeword_buf13[n*9+(16*C+3)],codeword_buf12[n*9+(16*C+3)],codeword_buf11[n*9+(16*C+3)],codeword_buf10[n*9+(16*C+3)],codeword_buf9[n*9+(16*C+3)],codeword_buf8[n*9+(16*C+3)],codeword_buf7[n*9+(16*C+3)],codeword_buf6[n*9+(16*C+3)],codeword_buf5[n*9+(16*C+3)],codeword_buf4[n*9+(16*C+3)],codeword_buf3[n*9+(16*C+3)],codeword_buf2[n*9+(16*C+3)],codeword_buf1[n*9+(16*C+3)],codeword_buf16[n*10+(16*C+3)],codeword_buf15[n*10+(16*C+3)],codeword_buf14[n*10+(16*C+3)],codeword_buf13[n*10+(16*C+3)],codeword_buf12[n*10+(16*C+3)],codeword_buf11[n*10+(16*C+3)],codeword_buf10[n*10+(16*C+3)],codeword_buf9[n*10+(16*C+3)],codeword_buf8[n*10+(16*C+3)],codeword_buf7[n*10+(16*C+3)],codeword_buf6[n*10+(16*C+3)],codeword_buf5[n*10+(16*C+3)],codeword_buf4[n*10+(16*C+3)],codeword_buf3[n*10+(16*C+3)],codeword_buf2[n*10+(16*C+3)],codeword_buf1[n*10+(16*C+3)],codeword_buf16[n*11+(16*C+3)],codeword_buf15[n*11+(16*C+3)],codeword_buf14[n*11+(16*C+3)],codeword_buf13[n*11+(16*C+3)],codeword_buf12[n*11+(16*C+3)],codeword_buf11[n*11+(16*C+3)],codeword_buf10[n*11+(16*C+3)],codeword_buf9[n*11+(16*C+3)],codeword_buf8[n*11+(16*C+3)],codeword_buf7[n*11+(16*C+3)],codeword_buf6[n*11+(16*C+3)],codeword_buf5[n*11+(16*C+3)],codeword_buf4[n*11+(16*C+3)],codeword_buf3[n*11+(16*C+3)],codeword_buf2[n*11+(16*C+3)],codeword_buf1[n*11+(16*C+3)],codeword_buf16[n*12+(16*C+3)],codeword_buf15[n*12+(16*C+3)],codeword_buf14[n*12+(16*C+3)],codeword_buf13[n*12+(16*C+3)],codeword_buf12[n*12+(16*C+3)],codeword_buf11[n*12+(16*C+3)],codeword_buf10[n*12+(16*C+3)],codeword_buf9[n*12+(16*C+3)],codeword_buf8[n*12+(16*C+3)],codeword_buf7[n*12+(16*C+3)],codeword_buf6[n*12+(16*C+3)],codeword_buf5[n*12+(16*C+3)],codeword_buf4[n*12+(16*C+3)],codeword_buf3[n*12+(16*C+3)],codeword_buf2[n*12+(16*C+3)],codeword_buf1[n*12+(16*C+3)],codeword_buf16[n*13+(16*C+3)],codeword_buf15[n*13+(16*C+3)],codeword_buf14[n*13+(16*C+3)],codeword_buf13[n*13+(16*C+3)],codeword_buf12[n*13+(16*C+3)],codeword_buf11[n*13+(16*C+3)],codeword_buf10[n*13+(16*C+3)],codeword_buf9[n*13+(16*C+3)],codeword_buf8[n*13+(16*C+3)],codeword_buf7[n*13+(16*C+3)],codeword_buf6[n*13+(16*C+3)],codeword_buf5[n*13+(16*C+3)],codeword_buf4[n*13+(16*C+3)],codeword_buf3[n*13+(16*C+3)],codeword_buf2[n*13+(16*C+3)],codeword_buf1[n*13+(16*C+3)],codeword_buf16[n*14+(16*C+3)],codeword_buf15[n*14+(16*C+3)],codeword_buf14[n*14+(16*C+3)],codeword_buf13[n*14+(16*C+3)],codeword_buf12[n*14+(16*C+3)],codeword_buf11[n*14+(16*C+3)],codeword_buf10[n*14+(16*C+3)],codeword_buf9[n*14+(16*C+3)],codeword_buf8[n*14+(16*C+3)],codeword_buf7[n*14+(16*C+3)],codeword_buf6[n*14+(16*C+3)],codeword_buf5[n*14+(16*C+3)],codeword_buf4[n*14+(16*C+3)],codeword_buf3[n*14+(16*C+3)],codeword_buf2[n*14+(16*C+3)],codeword_buf1[n*14+(16*C+3)],codeword_buf16[n*15+(16*C+3)],codeword_buf15[n*15+(16*C+3)],codeword_buf14[n*15+(16*C+3)],codeword_buf13[n*15+(16*C+3)],codeword_buf12[n*15+(16*C+3)],codeword_buf11[n*15+(16*C+3)],codeword_buf10[n*15+(16*C+3)],codeword_buf9[n*15+(16*C+3)],codeword_buf8[n*15+(16*C+3)],codeword_buf7[n*15+(16*C+3)],codeword_buf6[n*15+(16*C+3)],codeword_buf5[n*15+(16*C+3)],codeword_buf4[n*15+(16*C+3)],codeword_buf3[n*15+(16*C+3)],codeword_buf2[n*15+(16*C+3)],codeword_buf1[n*15+(16*C+3)]};
                            in_rec5 <= {codeword_buf16[n*0+(16*C+4)],codeword_buf15[n*0+(16*C+4)],codeword_buf14[n*0+(16*C+4)],codeword_buf13[n*0+(16*C+4)],codeword_buf12[n*0+(16*C+4)],codeword_buf11[n*0+(16*C+4)],codeword_buf10[n*0+(16*C+4)],codeword_buf9[n*0+(16*C+4)],codeword_buf8[n*0+(16*C+4)],codeword_buf7[n*0+(16*C+4)],codeword_buf6[n*0+(16*C+4)],codeword_buf5[n*0+(16*C+4)],codeword_buf4[n*0+(16*C+4)],codeword_buf3[n*0+(16*C+4)],codeword_buf2[n*0+(16*C+4)],codeword_buf1[n*0+(16*C+4)],codeword_buf16[n*1+(16*C+4)],codeword_buf15[n*1+(16*C+4)],codeword_buf14[n*1+(16*C+4)],codeword_buf13[n*1+(16*C+4)],codeword_buf12[n*1+(16*C+4)],codeword_buf11[n*1+(16*C+4)],codeword_buf10[n*1+(16*C+4)],codeword_buf9[n*1+(16*C+4)],codeword_buf8[n*1+(16*C+4)],codeword_buf7[n*1+(16*C+4)],codeword_buf6[n*1+(16*C+4)],codeword_buf5[n*1+(16*C+4)],codeword_buf4[n*1+(16*C+4)],codeword_buf3[n*1+(16*C+4)],codeword_buf2[n*1+(16*C+4)],codeword_buf1[n*1+(16*C+4)],codeword_buf16[n*2+(16*C+4)],codeword_buf15[n*2+(16*C+4)],codeword_buf14[n*2+(16*C+4)],codeword_buf13[n*2+(16*C+4)],codeword_buf12[n*2+(16*C+4)],codeword_buf11[n*2+(16*C+4)],codeword_buf10[n*2+(16*C+4)],codeword_buf9[n*2+(16*C+4)],codeword_buf8[n*2+(16*C+4)],codeword_buf7[n*2+(16*C+4)],codeword_buf6[n*2+(16*C+4)],codeword_buf5[n*2+(16*C+4)],codeword_buf4[n*2+(16*C+4)],codeword_buf3[n*2+(16*C+4)],codeword_buf2[n*2+(16*C+4)],codeword_buf1[n*2+(16*C+4)],codeword_buf16[n*3+(16*C+4)],codeword_buf15[n*3+(16*C+4)],codeword_buf14[n*3+(16*C+4)],codeword_buf13[n*3+(16*C+4)],codeword_buf12[n*3+(16*C+4)],codeword_buf11[n*3+(16*C+4)],codeword_buf10[n*3+(16*C+4)],codeword_buf9[n*3+(16*C+4)],codeword_buf8[n*3+(16*C+4)],codeword_buf7[n*3+(16*C+4)],codeword_buf6[n*3+(16*C+4)],codeword_buf5[n*3+(16*C+4)],codeword_buf4[n*3+(16*C+4)],codeword_buf3[n*3+(16*C+4)],codeword_buf2[n*3+(16*C+4)],codeword_buf1[n*3+(16*C+4)],codeword_buf16[n*4+(16*C+4)],codeword_buf15[n*4+(16*C+4)],codeword_buf14[n*4+(16*C+4)],codeword_buf13[n*4+(16*C+4)],codeword_buf12[n*4+(16*C+4)],codeword_buf11[n*4+(16*C+4)],codeword_buf10[n*4+(16*C+4)],codeword_buf9[n*4+(16*C+4)],codeword_buf8[n*4+(16*C+4)],codeword_buf7[n*4+(16*C+4)],codeword_buf6[n*4+(16*C+4)],codeword_buf5[n*4+(16*C+4)],codeword_buf4[n*4+(16*C+4)],codeword_buf3[n*4+(16*C+4)],codeword_buf2[n*4+(16*C+4)],codeword_buf1[n*4+(16*C+4)],codeword_buf16[n*5+(16*C+4)],codeword_buf15[n*5+(16*C+4)],codeword_buf14[n*5+(16*C+4)],codeword_buf13[n*5+(16*C+4)],codeword_buf12[n*5+(16*C+4)],codeword_buf11[n*5+(16*C+4)],codeword_buf10[n*5+(16*C+4)],codeword_buf9[n*5+(16*C+4)],codeword_buf8[n*5+(16*C+4)],codeword_buf7[n*5+(16*C+4)],codeword_buf6[n*5+(16*C+4)],codeword_buf5[n*5+(16*C+4)],codeword_buf4[n*5+(16*C+4)],codeword_buf3[n*5+(16*C+4)],codeword_buf2[n*5+(16*C+4)],codeword_buf1[n*5+(16*C+4)],codeword_buf16[n*6+(16*C+4)],codeword_buf15[n*6+(16*C+4)],codeword_buf14[n*6+(16*C+4)],codeword_buf13[n*6+(16*C+4)],codeword_buf12[n*6+(16*C+4)],codeword_buf11[n*6+(16*C+4)],codeword_buf10[n*6+(16*C+4)],codeword_buf9[n*6+(16*C+4)],codeword_buf8[n*6+(16*C+4)],codeword_buf7[n*6+(16*C+4)],codeword_buf6[n*6+(16*C+4)],codeword_buf5[n*6+(16*C+4)],codeword_buf4[n*6+(16*C+4)],codeword_buf3[n*6+(16*C+4)],codeword_buf2[n*6+(16*C+4)],codeword_buf1[n*6+(16*C+4)],codeword_buf16[n*7+(16*C+4)],codeword_buf15[n*7+(16*C+4)],codeword_buf14[n*7+(16*C+4)],codeword_buf13[n*7+(16*C+4)],codeword_buf12[n*7+(16*C+4)],codeword_buf11[n*7+(16*C+4)],codeword_buf10[n*7+(16*C+4)],codeword_buf9[n*7+(16*C+4)],codeword_buf8[n*7+(16*C+4)],codeword_buf7[n*7+(16*C+4)],codeword_buf6[n*7+(16*C+4)],codeword_buf5[n*7+(16*C+4)],codeword_buf4[n*7+(16*C+4)],codeword_buf3[n*7+(16*C+4)],codeword_buf2[n*7+(16*C+4)],codeword_buf1[n*7+(16*C+4)],codeword_buf16[n*8+(16*C+4)],codeword_buf15[n*8+(16*C+4)],codeword_buf14[n*8+(16*C+4)],codeword_buf13[n*8+(16*C+4)],codeword_buf12[n*8+(16*C+4)],codeword_buf11[n*8+(16*C+4)],codeword_buf10[n*8+(16*C+4)],codeword_buf9[n*8+(16*C+4)],codeword_buf8[n*8+(16*C+4)],codeword_buf7[n*8+(16*C+4)],codeword_buf6[n*8+(16*C+4)],codeword_buf5[n*8+(16*C+4)],codeword_buf4[n*8+(16*C+4)],codeword_buf3[n*8+(16*C+4)],codeword_buf2[n*8+(16*C+4)],codeword_buf1[n*8+(16*C+4)],codeword_buf16[n*9+(16*C+4)],codeword_buf15[n*9+(16*C+4)],codeword_buf14[n*9+(16*C+4)],codeword_buf13[n*9+(16*C+4)],codeword_buf12[n*9+(16*C+4)],codeword_buf11[n*9+(16*C+4)],codeword_buf10[n*9+(16*C+4)],codeword_buf9[n*9+(16*C+4)],codeword_buf8[n*9+(16*C+4)],codeword_buf7[n*9+(16*C+4)],codeword_buf6[n*9+(16*C+4)],codeword_buf5[n*9+(16*C+4)],codeword_buf4[n*9+(16*C+4)],codeword_buf3[n*9+(16*C+4)],codeword_buf2[n*9+(16*C+4)],codeword_buf1[n*9+(16*C+4)],codeword_buf16[n*10+(16*C+4)],codeword_buf15[n*10+(16*C+4)],codeword_buf14[n*10+(16*C+4)],codeword_buf13[n*10+(16*C+4)],codeword_buf12[n*10+(16*C+4)],codeword_buf11[n*10+(16*C+4)],codeword_buf10[n*10+(16*C+4)],codeword_buf9[n*10+(16*C+4)],codeword_buf8[n*10+(16*C+4)],codeword_buf7[n*10+(16*C+4)],codeword_buf6[n*10+(16*C+4)],codeword_buf5[n*10+(16*C+4)],codeword_buf4[n*10+(16*C+4)],codeword_buf3[n*10+(16*C+4)],codeword_buf2[n*10+(16*C+4)],codeword_buf1[n*10+(16*C+4)],codeword_buf16[n*11+(16*C+4)],codeword_buf15[n*11+(16*C+4)],codeword_buf14[n*11+(16*C+4)],codeword_buf13[n*11+(16*C+4)],codeword_buf12[n*11+(16*C+4)],codeword_buf11[n*11+(16*C+4)],codeword_buf10[n*11+(16*C+4)],codeword_buf9[n*11+(16*C+4)],codeword_buf8[n*11+(16*C+4)],codeword_buf7[n*11+(16*C+4)],codeword_buf6[n*11+(16*C+4)],codeword_buf5[n*11+(16*C+4)],codeword_buf4[n*11+(16*C+4)],codeword_buf3[n*11+(16*C+4)],codeword_buf2[n*11+(16*C+4)],codeword_buf1[n*11+(16*C+4)],codeword_buf16[n*12+(16*C+4)],codeword_buf15[n*12+(16*C+4)],codeword_buf14[n*12+(16*C+4)],codeword_buf13[n*12+(16*C+4)],codeword_buf12[n*12+(16*C+4)],codeword_buf11[n*12+(16*C+4)],codeword_buf10[n*12+(16*C+4)],codeword_buf9[n*12+(16*C+4)],codeword_buf8[n*12+(16*C+4)],codeword_buf7[n*12+(16*C+4)],codeword_buf6[n*12+(16*C+4)],codeword_buf5[n*12+(16*C+4)],codeword_buf4[n*12+(16*C+4)],codeword_buf3[n*12+(16*C+4)],codeword_buf2[n*12+(16*C+4)],codeword_buf1[n*12+(16*C+4)],codeword_buf16[n*13+(16*C+4)],codeword_buf15[n*13+(16*C+4)],codeword_buf14[n*13+(16*C+4)],codeword_buf13[n*13+(16*C+4)],codeword_buf12[n*13+(16*C+4)],codeword_buf11[n*13+(16*C+4)],codeword_buf10[n*13+(16*C+4)],codeword_buf9[n*13+(16*C+4)],codeword_buf8[n*13+(16*C+4)],codeword_buf7[n*13+(16*C+4)],codeword_buf6[n*13+(16*C+4)],codeword_buf5[n*13+(16*C+4)],codeword_buf4[n*13+(16*C+4)],codeword_buf3[n*13+(16*C+4)],codeword_buf2[n*13+(16*C+4)],codeword_buf1[n*13+(16*C+4)],codeword_buf16[n*14+(16*C+4)],codeword_buf15[n*14+(16*C+4)],codeword_buf14[n*14+(16*C+4)],codeword_buf13[n*14+(16*C+4)],codeword_buf12[n*14+(16*C+4)],codeword_buf11[n*14+(16*C+4)],codeword_buf10[n*14+(16*C+4)],codeword_buf9[n*14+(16*C+4)],codeword_buf8[n*14+(16*C+4)],codeword_buf7[n*14+(16*C+4)],codeword_buf6[n*14+(16*C+4)],codeword_buf5[n*14+(16*C+4)],codeword_buf4[n*14+(16*C+4)],codeword_buf3[n*14+(16*C+4)],codeword_buf2[n*14+(16*C+4)],codeword_buf1[n*14+(16*C+4)],codeword_buf16[n*15+(16*C+4)],codeword_buf15[n*15+(16*C+4)],codeword_buf14[n*15+(16*C+4)],codeword_buf13[n*15+(16*C+4)],codeword_buf12[n*15+(16*C+4)],codeword_buf11[n*15+(16*C+4)],codeword_buf10[n*15+(16*C+4)],codeword_buf9[n*15+(16*C+4)],codeword_buf8[n*15+(16*C+4)],codeword_buf7[n*15+(16*C+4)],codeword_buf6[n*15+(16*C+4)],codeword_buf5[n*15+(16*C+4)],codeword_buf4[n*15+(16*C+4)],codeword_buf3[n*15+(16*C+4)],codeword_buf2[n*15+(16*C+4)],codeword_buf1[n*15+(16*C+4)]};
                            in_rec6 <= {codeword_buf16[n*0+(16*C+5)],codeword_buf15[n*0+(16*C+5)],codeword_buf14[n*0+(16*C+5)],codeword_buf13[n*0+(16*C+5)],codeword_buf12[n*0+(16*C+5)],codeword_buf11[n*0+(16*C+5)],codeword_buf10[n*0+(16*C+5)],codeword_buf9[n*0+(16*C+5)],codeword_buf8[n*0+(16*C+5)],codeword_buf7[n*0+(16*C+5)],codeword_buf6[n*0+(16*C+5)],codeword_buf5[n*0+(16*C+5)],codeword_buf4[n*0+(16*C+5)],codeword_buf3[n*0+(16*C+5)],codeword_buf2[n*0+(16*C+5)],codeword_buf1[n*0+(16*C+5)],codeword_buf16[n*1+(16*C+5)],codeword_buf15[n*1+(16*C+5)],codeword_buf14[n*1+(16*C+5)],codeword_buf13[n*1+(16*C+5)],codeword_buf12[n*1+(16*C+5)],codeword_buf11[n*1+(16*C+5)],codeword_buf10[n*1+(16*C+5)],codeword_buf9[n*1+(16*C+5)],codeword_buf8[n*1+(16*C+5)],codeword_buf7[n*1+(16*C+5)],codeword_buf6[n*1+(16*C+5)],codeword_buf5[n*1+(16*C+5)],codeword_buf4[n*1+(16*C+5)],codeword_buf3[n*1+(16*C+5)],codeword_buf2[n*1+(16*C+5)],codeword_buf1[n*1+(16*C+5)],codeword_buf16[n*2+(16*C+5)],codeword_buf15[n*2+(16*C+5)],codeword_buf14[n*2+(16*C+5)],codeword_buf13[n*2+(16*C+5)],codeword_buf12[n*2+(16*C+5)],codeword_buf11[n*2+(16*C+5)],codeword_buf10[n*2+(16*C+5)],codeword_buf9[n*2+(16*C+5)],codeword_buf8[n*2+(16*C+5)],codeword_buf7[n*2+(16*C+5)],codeword_buf6[n*2+(16*C+5)],codeword_buf5[n*2+(16*C+5)],codeword_buf4[n*2+(16*C+5)],codeword_buf3[n*2+(16*C+5)],codeword_buf2[n*2+(16*C+5)],codeword_buf1[n*2+(16*C+5)],codeword_buf16[n*3+(16*C+5)],codeword_buf15[n*3+(16*C+5)],codeword_buf14[n*3+(16*C+5)],codeword_buf13[n*3+(16*C+5)],codeword_buf12[n*3+(16*C+5)],codeword_buf11[n*3+(16*C+5)],codeword_buf10[n*3+(16*C+5)],codeword_buf9[n*3+(16*C+5)],codeword_buf8[n*3+(16*C+5)],codeword_buf7[n*3+(16*C+5)],codeword_buf6[n*3+(16*C+5)],codeword_buf5[n*3+(16*C+5)],codeword_buf4[n*3+(16*C+5)],codeword_buf3[n*3+(16*C+5)],codeword_buf2[n*3+(16*C+5)],codeword_buf1[n*3+(16*C+5)],codeword_buf16[n*4+(16*C+5)],codeword_buf15[n*4+(16*C+5)],codeword_buf14[n*4+(16*C+5)],codeword_buf13[n*4+(16*C+5)],codeword_buf12[n*4+(16*C+5)],codeword_buf11[n*4+(16*C+5)],codeword_buf10[n*4+(16*C+5)],codeword_buf9[n*4+(16*C+5)],codeword_buf8[n*4+(16*C+5)],codeword_buf7[n*4+(16*C+5)],codeword_buf6[n*4+(16*C+5)],codeword_buf5[n*4+(16*C+5)],codeword_buf4[n*4+(16*C+5)],codeword_buf3[n*4+(16*C+5)],codeword_buf2[n*4+(16*C+5)],codeword_buf1[n*4+(16*C+5)],codeword_buf16[n*5+(16*C+5)],codeword_buf15[n*5+(16*C+5)],codeword_buf14[n*5+(16*C+5)],codeword_buf13[n*5+(16*C+5)],codeword_buf12[n*5+(16*C+5)],codeword_buf11[n*5+(16*C+5)],codeword_buf10[n*5+(16*C+5)],codeword_buf9[n*5+(16*C+5)],codeword_buf8[n*5+(16*C+5)],codeword_buf7[n*5+(16*C+5)],codeword_buf6[n*5+(16*C+5)],codeword_buf5[n*5+(16*C+5)],codeword_buf4[n*5+(16*C+5)],codeword_buf3[n*5+(16*C+5)],codeword_buf2[n*5+(16*C+5)],codeword_buf1[n*5+(16*C+5)],codeword_buf16[n*6+(16*C+5)],codeword_buf15[n*6+(16*C+5)],codeword_buf14[n*6+(16*C+5)],codeword_buf13[n*6+(16*C+5)],codeword_buf12[n*6+(16*C+5)],codeword_buf11[n*6+(16*C+5)],codeword_buf10[n*6+(16*C+5)],codeword_buf9[n*6+(16*C+5)],codeword_buf8[n*6+(16*C+5)],codeword_buf7[n*6+(16*C+5)],codeword_buf6[n*6+(16*C+5)],codeword_buf5[n*6+(16*C+5)],codeword_buf4[n*6+(16*C+5)],codeword_buf3[n*6+(16*C+5)],codeword_buf2[n*6+(16*C+5)],codeword_buf1[n*6+(16*C+5)],codeword_buf16[n*7+(16*C+5)],codeword_buf15[n*7+(16*C+5)],codeword_buf14[n*7+(16*C+5)],codeword_buf13[n*7+(16*C+5)],codeword_buf12[n*7+(16*C+5)],codeword_buf11[n*7+(16*C+5)],codeword_buf10[n*7+(16*C+5)],codeword_buf9[n*7+(16*C+5)],codeword_buf8[n*7+(16*C+5)],codeword_buf7[n*7+(16*C+5)],codeword_buf6[n*7+(16*C+5)],codeword_buf5[n*7+(16*C+5)],codeword_buf4[n*7+(16*C+5)],codeword_buf3[n*7+(16*C+5)],codeword_buf2[n*7+(16*C+5)],codeword_buf1[n*7+(16*C+5)],codeword_buf16[n*8+(16*C+5)],codeword_buf15[n*8+(16*C+5)],codeword_buf14[n*8+(16*C+5)],codeword_buf13[n*8+(16*C+5)],codeword_buf12[n*8+(16*C+5)],codeword_buf11[n*8+(16*C+5)],codeword_buf10[n*8+(16*C+5)],codeword_buf9[n*8+(16*C+5)],codeword_buf8[n*8+(16*C+5)],codeword_buf7[n*8+(16*C+5)],codeword_buf6[n*8+(16*C+5)],codeword_buf5[n*8+(16*C+5)],codeword_buf4[n*8+(16*C+5)],codeword_buf3[n*8+(16*C+5)],codeword_buf2[n*8+(16*C+5)],codeword_buf1[n*8+(16*C+5)],codeword_buf16[n*9+(16*C+5)],codeword_buf15[n*9+(16*C+5)],codeword_buf14[n*9+(16*C+5)],codeword_buf13[n*9+(16*C+5)],codeword_buf12[n*9+(16*C+5)],codeword_buf11[n*9+(16*C+5)],codeword_buf10[n*9+(16*C+5)],codeword_buf9[n*9+(16*C+5)],codeword_buf8[n*9+(16*C+5)],codeword_buf7[n*9+(16*C+5)],codeword_buf6[n*9+(16*C+5)],codeword_buf5[n*9+(16*C+5)],codeword_buf4[n*9+(16*C+5)],codeword_buf3[n*9+(16*C+5)],codeword_buf2[n*9+(16*C+5)],codeword_buf1[n*9+(16*C+5)],codeword_buf16[n*10+(16*C+5)],codeword_buf15[n*10+(16*C+5)],codeword_buf14[n*10+(16*C+5)],codeword_buf13[n*10+(16*C+5)],codeword_buf12[n*10+(16*C+5)],codeword_buf11[n*10+(16*C+5)],codeword_buf10[n*10+(16*C+5)],codeword_buf9[n*10+(16*C+5)],codeword_buf8[n*10+(16*C+5)],codeword_buf7[n*10+(16*C+5)],codeword_buf6[n*10+(16*C+5)],codeword_buf5[n*10+(16*C+5)],codeword_buf4[n*10+(16*C+5)],codeword_buf3[n*10+(16*C+5)],codeword_buf2[n*10+(16*C+5)],codeword_buf1[n*10+(16*C+5)],codeword_buf16[n*11+(16*C+5)],codeword_buf15[n*11+(16*C+5)],codeword_buf14[n*11+(16*C+5)],codeword_buf13[n*11+(16*C+5)],codeword_buf12[n*11+(16*C+5)],codeword_buf11[n*11+(16*C+5)],codeword_buf10[n*11+(16*C+5)],codeword_buf9[n*11+(16*C+5)],codeword_buf8[n*11+(16*C+5)],codeword_buf7[n*11+(16*C+5)],codeword_buf6[n*11+(16*C+5)],codeword_buf5[n*11+(16*C+5)],codeword_buf4[n*11+(16*C+5)],codeword_buf3[n*11+(16*C+5)],codeword_buf2[n*11+(16*C+5)],codeword_buf1[n*11+(16*C+5)],codeword_buf16[n*12+(16*C+5)],codeword_buf15[n*12+(16*C+5)],codeword_buf14[n*12+(16*C+5)],codeword_buf13[n*12+(16*C+5)],codeword_buf12[n*12+(16*C+5)],codeword_buf11[n*12+(16*C+5)],codeword_buf10[n*12+(16*C+5)],codeword_buf9[n*12+(16*C+5)],codeword_buf8[n*12+(16*C+5)],codeword_buf7[n*12+(16*C+5)],codeword_buf6[n*12+(16*C+5)],codeword_buf5[n*12+(16*C+5)],codeword_buf4[n*12+(16*C+5)],codeword_buf3[n*12+(16*C+5)],codeword_buf2[n*12+(16*C+5)],codeword_buf1[n*12+(16*C+5)],codeword_buf16[n*13+(16*C+5)],codeword_buf15[n*13+(16*C+5)],codeword_buf14[n*13+(16*C+5)],codeword_buf13[n*13+(16*C+5)],codeword_buf12[n*13+(16*C+5)],codeword_buf11[n*13+(16*C+5)],codeword_buf10[n*13+(16*C+5)],codeword_buf9[n*13+(16*C+5)],codeword_buf8[n*13+(16*C+5)],codeword_buf7[n*13+(16*C+5)],codeword_buf6[n*13+(16*C+5)],codeword_buf5[n*13+(16*C+5)],codeword_buf4[n*13+(16*C+5)],codeword_buf3[n*13+(16*C+5)],codeword_buf2[n*13+(16*C+5)],codeword_buf1[n*13+(16*C+5)],codeword_buf16[n*14+(16*C+5)],codeword_buf15[n*14+(16*C+5)],codeword_buf14[n*14+(16*C+5)],codeword_buf13[n*14+(16*C+5)],codeword_buf12[n*14+(16*C+5)],codeword_buf11[n*14+(16*C+5)],codeword_buf10[n*14+(16*C+5)],codeword_buf9[n*14+(16*C+5)],codeword_buf8[n*14+(16*C+5)],codeword_buf7[n*14+(16*C+5)],codeword_buf6[n*14+(16*C+5)],codeword_buf5[n*14+(16*C+5)],codeword_buf4[n*14+(16*C+5)],codeword_buf3[n*14+(16*C+5)],codeword_buf2[n*14+(16*C+5)],codeword_buf1[n*14+(16*C+5)],codeword_buf16[n*15+(16*C+5)],codeword_buf15[n*15+(16*C+5)],codeword_buf14[n*15+(16*C+5)],codeword_buf13[n*15+(16*C+5)],codeword_buf12[n*15+(16*C+5)],codeword_buf11[n*15+(16*C+5)],codeword_buf10[n*15+(16*C+5)],codeword_buf9[n*15+(16*C+5)],codeword_buf8[n*15+(16*C+5)],codeword_buf7[n*15+(16*C+5)],codeword_buf6[n*15+(16*C+5)],codeword_buf5[n*15+(16*C+5)],codeword_buf4[n*15+(16*C+5)],codeword_buf3[n*15+(16*C+5)],codeword_buf2[n*15+(16*C+5)],codeword_buf1[n*15+(16*C+5)]};
                            in_rec7 <= {codeword_buf16[n*0+(16*C+6)],codeword_buf15[n*0+(16*C+6)],codeword_buf14[n*0+(16*C+6)],codeword_buf13[n*0+(16*C+6)],codeword_buf12[n*0+(16*C+6)],codeword_buf11[n*0+(16*C+6)],codeword_buf10[n*0+(16*C+6)],codeword_buf9[n*0+(16*C+6)],codeword_buf8[n*0+(16*C+6)],codeword_buf7[n*0+(16*C+6)],codeword_buf6[n*0+(16*C+6)],codeword_buf5[n*0+(16*C+6)],codeword_buf4[n*0+(16*C+6)],codeword_buf3[n*0+(16*C+6)],codeword_buf2[n*0+(16*C+6)],codeword_buf1[n*0+(16*C+6)],codeword_buf16[n*1+(16*C+6)],codeword_buf15[n*1+(16*C+6)],codeword_buf14[n*1+(16*C+6)],codeword_buf13[n*1+(16*C+6)],codeword_buf12[n*1+(16*C+6)],codeword_buf11[n*1+(16*C+6)],codeword_buf10[n*1+(16*C+6)],codeword_buf9[n*1+(16*C+6)],codeword_buf8[n*1+(16*C+6)],codeword_buf7[n*1+(16*C+6)],codeword_buf6[n*1+(16*C+6)],codeword_buf5[n*1+(16*C+6)],codeword_buf4[n*1+(16*C+6)],codeword_buf3[n*1+(16*C+6)],codeword_buf2[n*1+(16*C+6)],codeword_buf1[n*1+(16*C+6)],codeword_buf16[n*2+(16*C+6)],codeword_buf15[n*2+(16*C+6)],codeword_buf14[n*2+(16*C+6)],codeword_buf13[n*2+(16*C+6)],codeword_buf12[n*2+(16*C+6)],codeword_buf11[n*2+(16*C+6)],codeword_buf10[n*2+(16*C+6)],codeword_buf9[n*2+(16*C+6)],codeword_buf8[n*2+(16*C+6)],codeword_buf7[n*2+(16*C+6)],codeword_buf6[n*2+(16*C+6)],codeword_buf5[n*2+(16*C+6)],codeword_buf4[n*2+(16*C+6)],codeword_buf3[n*2+(16*C+6)],codeword_buf2[n*2+(16*C+6)],codeword_buf1[n*2+(16*C+6)],codeword_buf16[n*3+(16*C+6)],codeword_buf15[n*3+(16*C+6)],codeword_buf14[n*3+(16*C+6)],codeword_buf13[n*3+(16*C+6)],codeword_buf12[n*3+(16*C+6)],codeword_buf11[n*3+(16*C+6)],codeword_buf10[n*3+(16*C+6)],codeword_buf9[n*3+(16*C+6)],codeword_buf8[n*3+(16*C+6)],codeword_buf7[n*3+(16*C+6)],codeword_buf6[n*3+(16*C+6)],codeword_buf5[n*3+(16*C+6)],codeword_buf4[n*3+(16*C+6)],codeword_buf3[n*3+(16*C+6)],codeword_buf2[n*3+(16*C+6)],codeword_buf1[n*3+(16*C+6)],codeword_buf16[n*4+(16*C+6)],codeword_buf15[n*4+(16*C+6)],codeword_buf14[n*4+(16*C+6)],codeword_buf13[n*4+(16*C+6)],codeword_buf12[n*4+(16*C+6)],codeword_buf11[n*4+(16*C+6)],codeword_buf10[n*4+(16*C+6)],codeword_buf9[n*4+(16*C+6)],codeword_buf8[n*4+(16*C+6)],codeword_buf7[n*4+(16*C+6)],codeword_buf6[n*4+(16*C+6)],codeword_buf5[n*4+(16*C+6)],codeword_buf4[n*4+(16*C+6)],codeword_buf3[n*4+(16*C+6)],codeword_buf2[n*4+(16*C+6)],codeword_buf1[n*4+(16*C+6)],codeword_buf16[n*5+(16*C+6)],codeword_buf15[n*5+(16*C+6)],codeword_buf14[n*5+(16*C+6)],codeword_buf13[n*5+(16*C+6)],codeword_buf12[n*5+(16*C+6)],codeword_buf11[n*5+(16*C+6)],codeword_buf10[n*5+(16*C+6)],codeword_buf9[n*5+(16*C+6)],codeword_buf8[n*5+(16*C+6)],codeword_buf7[n*5+(16*C+6)],codeword_buf6[n*5+(16*C+6)],codeword_buf5[n*5+(16*C+6)],codeword_buf4[n*5+(16*C+6)],codeword_buf3[n*5+(16*C+6)],codeword_buf2[n*5+(16*C+6)],codeword_buf1[n*5+(16*C+6)],codeword_buf16[n*6+(16*C+6)],codeword_buf15[n*6+(16*C+6)],codeword_buf14[n*6+(16*C+6)],codeword_buf13[n*6+(16*C+6)],codeword_buf12[n*6+(16*C+6)],codeword_buf11[n*6+(16*C+6)],codeword_buf10[n*6+(16*C+6)],codeword_buf9[n*6+(16*C+6)],codeword_buf8[n*6+(16*C+6)],codeword_buf7[n*6+(16*C+6)],codeword_buf6[n*6+(16*C+6)],codeword_buf5[n*6+(16*C+6)],codeword_buf4[n*6+(16*C+6)],codeword_buf3[n*6+(16*C+6)],codeword_buf2[n*6+(16*C+6)],codeword_buf1[n*6+(16*C+6)],codeword_buf16[n*7+(16*C+6)],codeword_buf15[n*7+(16*C+6)],codeword_buf14[n*7+(16*C+6)],codeword_buf13[n*7+(16*C+6)],codeword_buf12[n*7+(16*C+6)],codeword_buf11[n*7+(16*C+6)],codeword_buf10[n*7+(16*C+6)],codeword_buf9[n*7+(16*C+6)],codeword_buf8[n*7+(16*C+6)],codeword_buf7[n*7+(16*C+6)],codeword_buf6[n*7+(16*C+6)],codeword_buf5[n*7+(16*C+6)],codeword_buf4[n*7+(16*C+6)],codeword_buf3[n*7+(16*C+6)],codeword_buf2[n*7+(16*C+6)],codeword_buf1[n*7+(16*C+6)],codeword_buf16[n*8+(16*C+6)],codeword_buf15[n*8+(16*C+6)],codeword_buf14[n*8+(16*C+6)],codeword_buf13[n*8+(16*C+6)],codeword_buf12[n*8+(16*C+6)],codeword_buf11[n*8+(16*C+6)],codeword_buf10[n*8+(16*C+6)],codeword_buf9[n*8+(16*C+6)],codeword_buf8[n*8+(16*C+6)],codeword_buf7[n*8+(16*C+6)],codeword_buf6[n*8+(16*C+6)],codeword_buf5[n*8+(16*C+6)],codeword_buf4[n*8+(16*C+6)],codeword_buf3[n*8+(16*C+6)],codeword_buf2[n*8+(16*C+6)],codeword_buf1[n*8+(16*C+6)],codeword_buf16[n*9+(16*C+6)],codeword_buf15[n*9+(16*C+6)],codeword_buf14[n*9+(16*C+6)],codeword_buf13[n*9+(16*C+6)],codeword_buf12[n*9+(16*C+6)],codeword_buf11[n*9+(16*C+6)],codeword_buf10[n*9+(16*C+6)],codeword_buf9[n*9+(16*C+6)],codeword_buf8[n*9+(16*C+6)],codeword_buf7[n*9+(16*C+6)],codeword_buf6[n*9+(16*C+6)],codeword_buf5[n*9+(16*C+6)],codeword_buf4[n*9+(16*C+6)],codeword_buf3[n*9+(16*C+6)],codeword_buf2[n*9+(16*C+6)],codeword_buf1[n*9+(16*C+6)],codeword_buf16[n*10+(16*C+6)],codeword_buf15[n*10+(16*C+6)],codeword_buf14[n*10+(16*C+6)],codeword_buf13[n*10+(16*C+6)],codeword_buf12[n*10+(16*C+6)],codeword_buf11[n*10+(16*C+6)],codeword_buf10[n*10+(16*C+6)],codeword_buf9[n*10+(16*C+6)],codeword_buf8[n*10+(16*C+6)],codeword_buf7[n*10+(16*C+6)],codeword_buf6[n*10+(16*C+6)],codeword_buf5[n*10+(16*C+6)],codeword_buf4[n*10+(16*C+6)],codeword_buf3[n*10+(16*C+6)],codeword_buf2[n*10+(16*C+6)],codeword_buf1[n*10+(16*C+6)],codeword_buf16[n*11+(16*C+6)],codeword_buf15[n*11+(16*C+6)],codeword_buf14[n*11+(16*C+6)],codeword_buf13[n*11+(16*C+6)],codeword_buf12[n*11+(16*C+6)],codeword_buf11[n*11+(16*C+6)],codeword_buf10[n*11+(16*C+6)],codeword_buf9[n*11+(16*C+6)],codeword_buf8[n*11+(16*C+6)],codeword_buf7[n*11+(16*C+6)],codeword_buf6[n*11+(16*C+6)],codeword_buf5[n*11+(16*C+6)],codeword_buf4[n*11+(16*C+6)],codeword_buf3[n*11+(16*C+6)],codeword_buf2[n*11+(16*C+6)],codeword_buf1[n*11+(16*C+6)],codeword_buf16[n*12+(16*C+6)],codeword_buf15[n*12+(16*C+6)],codeword_buf14[n*12+(16*C+6)],codeword_buf13[n*12+(16*C+6)],codeword_buf12[n*12+(16*C+6)],codeword_buf11[n*12+(16*C+6)],codeword_buf10[n*12+(16*C+6)],codeword_buf9[n*12+(16*C+6)],codeword_buf8[n*12+(16*C+6)],codeword_buf7[n*12+(16*C+6)],codeword_buf6[n*12+(16*C+6)],codeword_buf5[n*12+(16*C+6)],codeword_buf4[n*12+(16*C+6)],codeword_buf3[n*12+(16*C+6)],codeword_buf2[n*12+(16*C+6)],codeword_buf1[n*12+(16*C+6)],codeword_buf16[n*13+(16*C+6)],codeword_buf15[n*13+(16*C+6)],codeword_buf14[n*13+(16*C+6)],codeword_buf13[n*13+(16*C+6)],codeword_buf12[n*13+(16*C+6)],codeword_buf11[n*13+(16*C+6)],codeword_buf10[n*13+(16*C+6)],codeword_buf9[n*13+(16*C+6)],codeword_buf8[n*13+(16*C+6)],codeword_buf7[n*13+(16*C+6)],codeword_buf6[n*13+(16*C+6)],codeword_buf5[n*13+(16*C+6)],codeword_buf4[n*13+(16*C+6)],codeword_buf3[n*13+(16*C+6)],codeword_buf2[n*13+(16*C+6)],codeword_buf1[n*13+(16*C+6)],codeword_buf16[n*14+(16*C+6)],codeword_buf15[n*14+(16*C+6)],codeword_buf14[n*14+(16*C+6)],codeword_buf13[n*14+(16*C+6)],codeword_buf12[n*14+(16*C+6)],codeword_buf11[n*14+(16*C+6)],codeword_buf10[n*14+(16*C+6)],codeword_buf9[n*14+(16*C+6)],codeword_buf8[n*14+(16*C+6)],codeword_buf7[n*14+(16*C+6)],codeword_buf6[n*14+(16*C+6)],codeword_buf5[n*14+(16*C+6)],codeword_buf4[n*14+(16*C+6)],codeword_buf3[n*14+(16*C+6)],codeword_buf2[n*14+(16*C+6)],codeword_buf1[n*14+(16*C+6)],codeword_buf16[n*15+(16*C+6)],codeword_buf15[n*15+(16*C+6)],codeword_buf14[n*15+(16*C+6)],codeword_buf13[n*15+(16*C+6)],codeword_buf12[n*15+(16*C+6)],codeword_buf11[n*15+(16*C+6)],codeword_buf10[n*15+(16*C+6)],codeword_buf9[n*15+(16*C+6)],codeword_buf8[n*15+(16*C+6)],codeword_buf7[n*15+(16*C+6)],codeword_buf6[n*15+(16*C+6)],codeword_buf5[n*15+(16*C+6)],codeword_buf4[n*15+(16*C+6)],codeword_buf3[n*15+(16*C+6)],codeword_buf2[n*15+(16*C+6)],codeword_buf1[n*15+(16*C+6)]};
                            in_rec8 <= {codeword_buf16[n*0+(16*C+7)],codeword_buf15[n*0+(16*C+7)],codeword_buf14[n*0+(16*C+7)],codeword_buf13[n*0+(16*C+7)],codeword_buf12[n*0+(16*C+7)],codeword_buf11[n*0+(16*C+7)],codeword_buf10[n*0+(16*C+7)],codeword_buf9[n*0+(16*C+7)],codeword_buf8[n*0+(16*C+7)],codeword_buf7[n*0+(16*C+7)],codeword_buf6[n*0+(16*C+7)],codeword_buf5[n*0+(16*C+7)],codeword_buf4[n*0+(16*C+7)],codeword_buf3[n*0+(16*C+7)],codeword_buf2[n*0+(16*C+7)],codeword_buf1[n*0+(16*C+7)],codeword_buf16[n*1+(16*C+7)],codeword_buf15[n*1+(16*C+7)],codeword_buf14[n*1+(16*C+7)],codeword_buf13[n*1+(16*C+7)],codeword_buf12[n*1+(16*C+7)],codeword_buf11[n*1+(16*C+7)],codeword_buf10[n*1+(16*C+7)],codeword_buf9[n*1+(16*C+7)],codeword_buf8[n*1+(16*C+7)],codeword_buf7[n*1+(16*C+7)],codeword_buf6[n*1+(16*C+7)],codeword_buf5[n*1+(16*C+7)],codeword_buf4[n*1+(16*C+7)],codeword_buf3[n*1+(16*C+7)],codeword_buf2[n*1+(16*C+7)],codeword_buf1[n*1+(16*C+7)],codeword_buf16[n*2+(16*C+7)],codeword_buf15[n*2+(16*C+7)],codeword_buf14[n*2+(16*C+7)],codeword_buf13[n*2+(16*C+7)],codeword_buf12[n*2+(16*C+7)],codeword_buf11[n*2+(16*C+7)],codeword_buf10[n*2+(16*C+7)],codeword_buf9[n*2+(16*C+7)],codeword_buf8[n*2+(16*C+7)],codeword_buf7[n*2+(16*C+7)],codeword_buf6[n*2+(16*C+7)],codeword_buf5[n*2+(16*C+7)],codeword_buf4[n*2+(16*C+7)],codeword_buf3[n*2+(16*C+7)],codeword_buf2[n*2+(16*C+7)],codeword_buf1[n*2+(16*C+7)],codeword_buf16[n*3+(16*C+7)],codeword_buf15[n*3+(16*C+7)],codeword_buf14[n*3+(16*C+7)],codeword_buf13[n*3+(16*C+7)],codeword_buf12[n*3+(16*C+7)],codeword_buf11[n*3+(16*C+7)],codeword_buf10[n*3+(16*C+7)],codeword_buf9[n*3+(16*C+7)],codeword_buf8[n*3+(16*C+7)],codeword_buf7[n*3+(16*C+7)],codeword_buf6[n*3+(16*C+7)],codeword_buf5[n*3+(16*C+7)],codeword_buf4[n*3+(16*C+7)],codeword_buf3[n*3+(16*C+7)],codeword_buf2[n*3+(16*C+7)],codeword_buf1[n*3+(16*C+7)],codeword_buf16[n*4+(16*C+7)],codeword_buf15[n*4+(16*C+7)],codeword_buf14[n*4+(16*C+7)],codeword_buf13[n*4+(16*C+7)],codeword_buf12[n*4+(16*C+7)],codeword_buf11[n*4+(16*C+7)],codeword_buf10[n*4+(16*C+7)],codeword_buf9[n*4+(16*C+7)],codeword_buf8[n*4+(16*C+7)],codeword_buf7[n*4+(16*C+7)],codeword_buf6[n*4+(16*C+7)],codeword_buf5[n*4+(16*C+7)],codeword_buf4[n*4+(16*C+7)],codeword_buf3[n*4+(16*C+7)],codeword_buf2[n*4+(16*C+7)],codeword_buf1[n*4+(16*C+7)],codeword_buf16[n*5+(16*C+7)],codeword_buf15[n*5+(16*C+7)],codeword_buf14[n*5+(16*C+7)],codeword_buf13[n*5+(16*C+7)],codeword_buf12[n*5+(16*C+7)],codeword_buf11[n*5+(16*C+7)],codeword_buf10[n*5+(16*C+7)],codeword_buf9[n*5+(16*C+7)],codeword_buf8[n*5+(16*C+7)],codeword_buf7[n*5+(16*C+7)],codeword_buf6[n*5+(16*C+7)],codeword_buf5[n*5+(16*C+7)],codeword_buf4[n*5+(16*C+7)],codeword_buf3[n*5+(16*C+7)],codeword_buf2[n*5+(16*C+7)],codeword_buf1[n*5+(16*C+7)],codeword_buf16[n*6+(16*C+7)],codeword_buf15[n*6+(16*C+7)],codeword_buf14[n*6+(16*C+7)],codeword_buf13[n*6+(16*C+7)],codeword_buf12[n*6+(16*C+7)],codeword_buf11[n*6+(16*C+7)],codeword_buf10[n*6+(16*C+7)],codeword_buf9[n*6+(16*C+7)],codeword_buf8[n*6+(16*C+7)],codeword_buf7[n*6+(16*C+7)],codeword_buf6[n*6+(16*C+7)],codeword_buf5[n*6+(16*C+7)],codeword_buf4[n*6+(16*C+7)],codeword_buf3[n*6+(16*C+7)],codeword_buf2[n*6+(16*C+7)],codeword_buf1[n*6+(16*C+7)],codeword_buf16[n*7+(16*C+7)],codeword_buf15[n*7+(16*C+7)],codeword_buf14[n*7+(16*C+7)],codeword_buf13[n*7+(16*C+7)],codeword_buf12[n*7+(16*C+7)],codeword_buf11[n*7+(16*C+7)],codeword_buf10[n*7+(16*C+7)],codeword_buf9[n*7+(16*C+7)],codeword_buf8[n*7+(16*C+7)],codeword_buf7[n*7+(16*C+7)],codeword_buf6[n*7+(16*C+7)],codeword_buf5[n*7+(16*C+7)],codeword_buf4[n*7+(16*C+7)],codeword_buf3[n*7+(16*C+7)],codeword_buf2[n*7+(16*C+7)],codeword_buf1[n*7+(16*C+7)],codeword_buf16[n*8+(16*C+7)],codeword_buf15[n*8+(16*C+7)],codeword_buf14[n*8+(16*C+7)],codeword_buf13[n*8+(16*C+7)],codeword_buf12[n*8+(16*C+7)],codeword_buf11[n*8+(16*C+7)],codeword_buf10[n*8+(16*C+7)],codeword_buf9[n*8+(16*C+7)],codeword_buf8[n*8+(16*C+7)],codeword_buf7[n*8+(16*C+7)],codeword_buf6[n*8+(16*C+7)],codeword_buf5[n*8+(16*C+7)],codeword_buf4[n*8+(16*C+7)],codeword_buf3[n*8+(16*C+7)],codeword_buf2[n*8+(16*C+7)],codeword_buf1[n*8+(16*C+7)],codeword_buf16[n*9+(16*C+7)],codeword_buf15[n*9+(16*C+7)],codeword_buf14[n*9+(16*C+7)],codeword_buf13[n*9+(16*C+7)],codeword_buf12[n*9+(16*C+7)],codeword_buf11[n*9+(16*C+7)],codeword_buf10[n*9+(16*C+7)],codeword_buf9[n*9+(16*C+7)],codeword_buf8[n*9+(16*C+7)],codeword_buf7[n*9+(16*C+7)],codeword_buf6[n*9+(16*C+7)],codeword_buf5[n*9+(16*C+7)],codeword_buf4[n*9+(16*C+7)],codeword_buf3[n*9+(16*C+7)],codeword_buf2[n*9+(16*C+7)],codeword_buf1[n*9+(16*C+7)],codeword_buf16[n*10+(16*C+7)],codeword_buf15[n*10+(16*C+7)],codeword_buf14[n*10+(16*C+7)],codeword_buf13[n*10+(16*C+7)],codeword_buf12[n*10+(16*C+7)],codeword_buf11[n*10+(16*C+7)],codeword_buf10[n*10+(16*C+7)],codeword_buf9[n*10+(16*C+7)],codeword_buf8[n*10+(16*C+7)],codeword_buf7[n*10+(16*C+7)],codeword_buf6[n*10+(16*C+7)],codeword_buf5[n*10+(16*C+7)],codeword_buf4[n*10+(16*C+7)],codeword_buf3[n*10+(16*C+7)],codeword_buf2[n*10+(16*C+7)],codeword_buf1[n*10+(16*C+7)],codeword_buf16[n*11+(16*C+7)],codeword_buf15[n*11+(16*C+7)],codeword_buf14[n*11+(16*C+7)],codeword_buf13[n*11+(16*C+7)],codeword_buf12[n*11+(16*C+7)],codeword_buf11[n*11+(16*C+7)],codeword_buf10[n*11+(16*C+7)],codeword_buf9[n*11+(16*C+7)],codeword_buf8[n*11+(16*C+7)],codeword_buf7[n*11+(16*C+7)],codeword_buf6[n*11+(16*C+7)],codeword_buf5[n*11+(16*C+7)],codeword_buf4[n*11+(16*C+7)],codeword_buf3[n*11+(16*C+7)],codeword_buf2[n*11+(16*C+7)],codeword_buf1[n*11+(16*C+7)],codeword_buf16[n*12+(16*C+7)],codeword_buf15[n*12+(16*C+7)],codeword_buf14[n*12+(16*C+7)],codeword_buf13[n*12+(16*C+7)],codeword_buf12[n*12+(16*C+7)],codeword_buf11[n*12+(16*C+7)],codeword_buf10[n*12+(16*C+7)],codeword_buf9[n*12+(16*C+7)],codeword_buf8[n*12+(16*C+7)],codeword_buf7[n*12+(16*C+7)],codeword_buf6[n*12+(16*C+7)],codeword_buf5[n*12+(16*C+7)],codeword_buf4[n*12+(16*C+7)],codeword_buf3[n*12+(16*C+7)],codeword_buf2[n*12+(16*C+7)],codeword_buf1[n*12+(16*C+7)],codeword_buf16[n*13+(16*C+7)],codeword_buf15[n*13+(16*C+7)],codeword_buf14[n*13+(16*C+7)],codeword_buf13[n*13+(16*C+7)],codeword_buf12[n*13+(16*C+7)],codeword_buf11[n*13+(16*C+7)],codeword_buf10[n*13+(16*C+7)],codeword_buf9[n*13+(16*C+7)],codeword_buf8[n*13+(16*C+7)],codeword_buf7[n*13+(16*C+7)],codeword_buf6[n*13+(16*C+7)],codeword_buf5[n*13+(16*C+7)],codeword_buf4[n*13+(16*C+7)],codeword_buf3[n*13+(16*C+7)],codeword_buf2[n*13+(16*C+7)],codeword_buf1[n*13+(16*C+7)],codeword_buf16[n*14+(16*C+7)],codeword_buf15[n*14+(16*C+7)],codeword_buf14[n*14+(16*C+7)],codeword_buf13[n*14+(16*C+7)],codeword_buf12[n*14+(16*C+7)],codeword_buf11[n*14+(16*C+7)],codeword_buf10[n*14+(16*C+7)],codeword_buf9[n*14+(16*C+7)],codeword_buf8[n*14+(16*C+7)],codeword_buf7[n*14+(16*C+7)],codeword_buf6[n*14+(16*C+7)],codeword_buf5[n*14+(16*C+7)],codeword_buf4[n*14+(16*C+7)],codeword_buf3[n*14+(16*C+7)],codeword_buf2[n*14+(16*C+7)],codeword_buf1[n*14+(16*C+7)],codeword_buf16[n*15+(16*C+7)],codeword_buf15[n*15+(16*C+7)],codeword_buf14[n*15+(16*C+7)],codeword_buf13[n*15+(16*C+7)],codeword_buf12[n*15+(16*C+7)],codeword_buf11[n*15+(16*C+7)],codeword_buf10[n*15+(16*C+7)],codeword_buf9[n*15+(16*C+7)],codeword_buf8[n*15+(16*C+7)],codeword_buf7[n*15+(16*C+7)],codeword_buf6[n*15+(16*C+7)],codeword_buf5[n*15+(16*C+7)],codeword_buf4[n*15+(16*C+7)],codeword_buf3[n*15+(16*C+7)],codeword_buf2[n*15+(16*C+7)],codeword_buf1[n*15+(16*C+7)]};
                            in_rec9 <= {codeword_buf16[n*0+(16*C+8)],codeword_buf15[n*0+(16*C+8)],codeword_buf14[n*0+(16*C+8)],codeword_buf13[n*0+(16*C+8)],codeword_buf12[n*0+(16*C+8)],codeword_buf11[n*0+(16*C+8)],codeword_buf10[n*0+(16*C+8)],codeword_buf9[n*0+(16*C+8)],codeword_buf8[n*0+(16*C+8)],codeword_buf7[n*0+(16*C+8)],codeword_buf6[n*0+(16*C+8)],codeword_buf5[n*0+(16*C+8)],codeword_buf4[n*0+(16*C+8)],codeword_buf3[n*0+(16*C+8)],codeword_buf2[n*0+(16*C+8)],codeword_buf1[n*0+(16*C+8)],codeword_buf16[n*1+(16*C+8)],codeword_buf15[n*1+(16*C+8)],codeword_buf14[n*1+(16*C+8)],codeword_buf13[n*1+(16*C+8)],codeword_buf12[n*1+(16*C+8)],codeword_buf11[n*1+(16*C+8)],codeword_buf10[n*1+(16*C+8)],codeword_buf9[n*1+(16*C+8)],codeword_buf8[n*1+(16*C+8)],codeword_buf7[n*1+(16*C+8)],codeword_buf6[n*1+(16*C+8)],codeword_buf5[n*1+(16*C+8)],codeword_buf4[n*1+(16*C+8)],codeword_buf3[n*1+(16*C+8)],codeword_buf2[n*1+(16*C+8)],codeword_buf1[n*1+(16*C+8)],codeword_buf16[n*2+(16*C+8)],codeword_buf15[n*2+(16*C+8)],codeword_buf14[n*2+(16*C+8)],codeword_buf13[n*2+(16*C+8)],codeword_buf12[n*2+(16*C+8)],codeword_buf11[n*2+(16*C+8)],codeword_buf10[n*2+(16*C+8)],codeword_buf9[n*2+(16*C+8)],codeword_buf8[n*2+(16*C+8)],codeword_buf7[n*2+(16*C+8)],codeword_buf6[n*2+(16*C+8)],codeword_buf5[n*2+(16*C+8)],codeword_buf4[n*2+(16*C+8)],codeword_buf3[n*2+(16*C+8)],codeword_buf2[n*2+(16*C+8)],codeword_buf1[n*2+(16*C+8)],codeword_buf16[n*3+(16*C+8)],codeword_buf15[n*3+(16*C+8)],codeword_buf14[n*3+(16*C+8)],codeword_buf13[n*3+(16*C+8)],codeword_buf12[n*3+(16*C+8)],codeword_buf11[n*3+(16*C+8)],codeword_buf10[n*3+(16*C+8)],codeword_buf9[n*3+(16*C+8)],codeword_buf8[n*3+(16*C+8)],codeword_buf7[n*3+(16*C+8)],codeword_buf6[n*3+(16*C+8)],codeword_buf5[n*3+(16*C+8)],codeword_buf4[n*3+(16*C+8)],codeword_buf3[n*3+(16*C+8)],codeword_buf2[n*3+(16*C+8)],codeword_buf1[n*3+(16*C+8)],codeword_buf16[n*4+(16*C+8)],codeword_buf15[n*4+(16*C+8)],codeword_buf14[n*4+(16*C+8)],codeword_buf13[n*4+(16*C+8)],codeword_buf12[n*4+(16*C+8)],codeword_buf11[n*4+(16*C+8)],codeword_buf10[n*4+(16*C+8)],codeword_buf9[n*4+(16*C+8)],codeword_buf8[n*4+(16*C+8)],codeword_buf7[n*4+(16*C+8)],codeword_buf6[n*4+(16*C+8)],codeword_buf5[n*4+(16*C+8)],codeword_buf4[n*4+(16*C+8)],codeword_buf3[n*4+(16*C+8)],codeword_buf2[n*4+(16*C+8)],codeword_buf1[n*4+(16*C+8)],codeword_buf16[n*5+(16*C+8)],codeword_buf15[n*5+(16*C+8)],codeword_buf14[n*5+(16*C+8)],codeword_buf13[n*5+(16*C+8)],codeword_buf12[n*5+(16*C+8)],codeword_buf11[n*5+(16*C+8)],codeword_buf10[n*5+(16*C+8)],codeword_buf9[n*5+(16*C+8)],codeword_buf8[n*5+(16*C+8)],codeword_buf7[n*5+(16*C+8)],codeword_buf6[n*5+(16*C+8)],codeword_buf5[n*5+(16*C+8)],codeword_buf4[n*5+(16*C+8)],codeword_buf3[n*5+(16*C+8)],codeword_buf2[n*5+(16*C+8)],codeword_buf1[n*5+(16*C+8)],codeword_buf16[n*6+(16*C+8)],codeword_buf15[n*6+(16*C+8)],codeword_buf14[n*6+(16*C+8)],codeword_buf13[n*6+(16*C+8)],codeword_buf12[n*6+(16*C+8)],codeword_buf11[n*6+(16*C+8)],codeword_buf10[n*6+(16*C+8)],codeword_buf9[n*6+(16*C+8)],codeword_buf8[n*6+(16*C+8)],codeword_buf7[n*6+(16*C+8)],codeword_buf6[n*6+(16*C+8)],codeword_buf5[n*6+(16*C+8)],codeword_buf4[n*6+(16*C+8)],codeword_buf3[n*6+(16*C+8)],codeword_buf2[n*6+(16*C+8)],codeword_buf1[n*6+(16*C+8)],codeword_buf16[n*7+(16*C+8)],codeword_buf15[n*7+(16*C+8)],codeword_buf14[n*7+(16*C+8)],codeword_buf13[n*7+(16*C+8)],codeword_buf12[n*7+(16*C+8)],codeword_buf11[n*7+(16*C+8)],codeword_buf10[n*7+(16*C+8)],codeword_buf9[n*7+(16*C+8)],codeword_buf8[n*7+(16*C+8)],codeword_buf7[n*7+(16*C+8)],codeword_buf6[n*7+(16*C+8)],codeword_buf5[n*7+(16*C+8)],codeword_buf4[n*7+(16*C+8)],codeword_buf3[n*7+(16*C+8)],codeword_buf2[n*7+(16*C+8)],codeword_buf1[n*7+(16*C+8)],codeword_buf16[n*8+(16*C+8)],codeword_buf15[n*8+(16*C+8)],codeword_buf14[n*8+(16*C+8)],codeword_buf13[n*8+(16*C+8)],codeword_buf12[n*8+(16*C+8)],codeword_buf11[n*8+(16*C+8)],codeword_buf10[n*8+(16*C+8)],codeword_buf9[n*8+(16*C+8)],codeword_buf8[n*8+(16*C+8)],codeword_buf7[n*8+(16*C+8)],codeword_buf6[n*8+(16*C+8)],codeword_buf5[n*8+(16*C+8)],codeword_buf4[n*8+(16*C+8)],codeword_buf3[n*8+(16*C+8)],codeword_buf2[n*8+(16*C+8)],codeword_buf1[n*8+(16*C+8)],codeword_buf16[n*9+(16*C+8)],codeword_buf15[n*9+(16*C+8)],codeword_buf14[n*9+(16*C+8)],codeword_buf13[n*9+(16*C+8)],codeword_buf12[n*9+(16*C+8)],codeword_buf11[n*9+(16*C+8)],codeword_buf10[n*9+(16*C+8)],codeword_buf9[n*9+(16*C+8)],codeword_buf8[n*9+(16*C+8)],codeword_buf7[n*9+(16*C+8)],codeword_buf6[n*9+(16*C+8)],codeword_buf5[n*9+(16*C+8)],codeword_buf4[n*9+(16*C+8)],codeword_buf3[n*9+(16*C+8)],codeword_buf2[n*9+(16*C+8)],codeword_buf1[n*9+(16*C+8)],codeword_buf16[n*10+(16*C+8)],codeword_buf15[n*10+(16*C+8)],codeword_buf14[n*10+(16*C+8)],codeword_buf13[n*10+(16*C+8)],codeword_buf12[n*10+(16*C+8)],codeword_buf11[n*10+(16*C+8)],codeword_buf10[n*10+(16*C+8)],codeword_buf9[n*10+(16*C+8)],codeword_buf8[n*10+(16*C+8)],codeword_buf7[n*10+(16*C+8)],codeword_buf6[n*10+(16*C+8)],codeword_buf5[n*10+(16*C+8)],codeword_buf4[n*10+(16*C+8)],codeword_buf3[n*10+(16*C+8)],codeword_buf2[n*10+(16*C+8)],codeword_buf1[n*10+(16*C+8)],codeword_buf16[n*11+(16*C+8)],codeword_buf15[n*11+(16*C+8)],codeword_buf14[n*11+(16*C+8)],codeword_buf13[n*11+(16*C+8)],codeword_buf12[n*11+(16*C+8)],codeword_buf11[n*11+(16*C+8)],codeword_buf10[n*11+(16*C+8)],codeword_buf9[n*11+(16*C+8)],codeword_buf8[n*11+(16*C+8)],codeword_buf7[n*11+(16*C+8)],codeword_buf6[n*11+(16*C+8)],codeword_buf5[n*11+(16*C+8)],codeword_buf4[n*11+(16*C+8)],codeword_buf3[n*11+(16*C+8)],codeword_buf2[n*11+(16*C+8)],codeword_buf1[n*11+(16*C+8)],codeword_buf16[n*12+(16*C+8)],codeword_buf15[n*12+(16*C+8)],codeword_buf14[n*12+(16*C+8)],codeword_buf13[n*12+(16*C+8)],codeword_buf12[n*12+(16*C+8)],codeword_buf11[n*12+(16*C+8)],codeword_buf10[n*12+(16*C+8)],codeword_buf9[n*12+(16*C+8)],codeword_buf8[n*12+(16*C+8)],codeword_buf7[n*12+(16*C+8)],codeword_buf6[n*12+(16*C+8)],codeword_buf5[n*12+(16*C+8)],codeword_buf4[n*12+(16*C+8)],codeword_buf3[n*12+(16*C+8)],codeword_buf2[n*12+(16*C+8)],codeword_buf1[n*12+(16*C+8)],codeword_buf16[n*13+(16*C+8)],codeword_buf15[n*13+(16*C+8)],codeword_buf14[n*13+(16*C+8)],codeword_buf13[n*13+(16*C+8)],codeword_buf12[n*13+(16*C+8)],codeword_buf11[n*13+(16*C+8)],codeword_buf10[n*13+(16*C+8)],codeword_buf9[n*13+(16*C+8)],codeword_buf8[n*13+(16*C+8)],codeword_buf7[n*13+(16*C+8)],codeword_buf6[n*13+(16*C+8)],codeword_buf5[n*13+(16*C+8)],codeword_buf4[n*13+(16*C+8)],codeword_buf3[n*13+(16*C+8)],codeword_buf2[n*13+(16*C+8)],codeword_buf1[n*13+(16*C+8)],codeword_buf16[n*14+(16*C+8)],codeword_buf15[n*14+(16*C+8)],codeword_buf14[n*14+(16*C+8)],codeword_buf13[n*14+(16*C+8)],codeword_buf12[n*14+(16*C+8)],codeword_buf11[n*14+(16*C+8)],codeword_buf10[n*14+(16*C+8)],codeword_buf9[n*14+(16*C+8)],codeword_buf8[n*14+(16*C+8)],codeword_buf7[n*14+(16*C+8)],codeword_buf6[n*14+(16*C+8)],codeword_buf5[n*14+(16*C+8)],codeword_buf4[n*14+(16*C+8)],codeword_buf3[n*14+(16*C+8)],codeword_buf2[n*14+(16*C+8)],codeword_buf1[n*14+(16*C+8)],codeword_buf16[n*15+(16*C+8)],codeword_buf15[n*15+(16*C+8)],codeword_buf14[n*15+(16*C+8)],codeword_buf13[n*15+(16*C+8)],codeword_buf12[n*15+(16*C+8)],codeword_buf11[n*15+(16*C+8)],codeword_buf10[n*15+(16*C+8)],codeword_buf9[n*15+(16*C+8)],codeword_buf8[n*15+(16*C+8)],codeword_buf7[n*15+(16*C+8)],codeword_buf6[n*15+(16*C+8)],codeword_buf5[n*15+(16*C+8)],codeword_buf4[n*15+(16*C+8)],codeword_buf3[n*15+(16*C+8)],codeword_buf2[n*15+(16*C+8)],codeword_buf1[n*15+(16*C+8)]};
                            in_rec10 <= {codeword_buf16[n*0+(16*C+9)],codeword_buf15[n*0+(16*C+9)],codeword_buf14[n*0+(16*C+9)],codeword_buf13[n*0+(16*C+9)],codeword_buf12[n*0+(16*C+9)],codeword_buf11[n*0+(16*C+9)],codeword_buf10[n*0+(16*C+9)],codeword_buf9[n*0+(16*C+9)],codeword_buf8[n*0+(16*C+9)],codeword_buf7[n*0+(16*C+9)],codeword_buf6[n*0+(16*C+9)],codeword_buf5[n*0+(16*C+9)],codeword_buf4[n*0+(16*C+9)],codeword_buf3[n*0+(16*C+9)],codeword_buf2[n*0+(16*C+9)],codeword_buf1[n*0+(16*C+9)],codeword_buf16[n*1+(16*C+9)],codeword_buf15[n*1+(16*C+9)],codeword_buf14[n*1+(16*C+9)],codeword_buf13[n*1+(16*C+9)],codeword_buf12[n*1+(16*C+9)],codeword_buf11[n*1+(16*C+9)],codeword_buf10[n*1+(16*C+9)],codeword_buf9[n*1+(16*C+9)],codeword_buf8[n*1+(16*C+9)],codeword_buf7[n*1+(16*C+9)],codeword_buf6[n*1+(16*C+9)],codeword_buf5[n*1+(16*C+9)],codeword_buf4[n*1+(16*C+9)],codeword_buf3[n*1+(16*C+9)],codeword_buf2[n*1+(16*C+9)],codeword_buf1[n*1+(16*C+9)],codeword_buf16[n*2+(16*C+9)],codeword_buf15[n*2+(16*C+9)],codeword_buf14[n*2+(16*C+9)],codeword_buf13[n*2+(16*C+9)],codeword_buf12[n*2+(16*C+9)],codeword_buf11[n*2+(16*C+9)],codeword_buf10[n*2+(16*C+9)],codeword_buf9[n*2+(16*C+9)],codeword_buf8[n*2+(16*C+9)],codeword_buf7[n*2+(16*C+9)],codeword_buf6[n*2+(16*C+9)],codeword_buf5[n*2+(16*C+9)],codeword_buf4[n*2+(16*C+9)],codeword_buf3[n*2+(16*C+9)],codeword_buf2[n*2+(16*C+9)],codeword_buf1[n*2+(16*C+9)],codeword_buf16[n*3+(16*C+9)],codeword_buf15[n*3+(16*C+9)],codeword_buf14[n*3+(16*C+9)],codeword_buf13[n*3+(16*C+9)],codeword_buf12[n*3+(16*C+9)],codeword_buf11[n*3+(16*C+9)],codeword_buf10[n*3+(16*C+9)],codeword_buf9[n*3+(16*C+9)],codeword_buf8[n*3+(16*C+9)],codeword_buf7[n*3+(16*C+9)],codeword_buf6[n*3+(16*C+9)],codeword_buf5[n*3+(16*C+9)],codeword_buf4[n*3+(16*C+9)],codeword_buf3[n*3+(16*C+9)],codeword_buf2[n*3+(16*C+9)],codeword_buf1[n*3+(16*C+9)],codeword_buf16[n*4+(16*C+9)],codeword_buf15[n*4+(16*C+9)],codeword_buf14[n*4+(16*C+9)],codeword_buf13[n*4+(16*C+9)],codeword_buf12[n*4+(16*C+9)],codeword_buf11[n*4+(16*C+9)],codeword_buf10[n*4+(16*C+9)],codeword_buf9[n*4+(16*C+9)],codeword_buf8[n*4+(16*C+9)],codeword_buf7[n*4+(16*C+9)],codeword_buf6[n*4+(16*C+9)],codeword_buf5[n*4+(16*C+9)],codeword_buf4[n*4+(16*C+9)],codeword_buf3[n*4+(16*C+9)],codeword_buf2[n*4+(16*C+9)],codeword_buf1[n*4+(16*C+9)],codeword_buf16[n*5+(16*C+9)],codeword_buf15[n*5+(16*C+9)],codeword_buf14[n*5+(16*C+9)],codeword_buf13[n*5+(16*C+9)],codeword_buf12[n*5+(16*C+9)],codeword_buf11[n*5+(16*C+9)],codeword_buf10[n*5+(16*C+9)],codeword_buf9[n*5+(16*C+9)],codeword_buf8[n*5+(16*C+9)],codeword_buf7[n*5+(16*C+9)],codeword_buf6[n*5+(16*C+9)],codeword_buf5[n*5+(16*C+9)],codeword_buf4[n*5+(16*C+9)],codeword_buf3[n*5+(16*C+9)],codeword_buf2[n*5+(16*C+9)],codeword_buf1[n*5+(16*C+9)],codeword_buf16[n*6+(16*C+9)],codeword_buf15[n*6+(16*C+9)],codeword_buf14[n*6+(16*C+9)],codeword_buf13[n*6+(16*C+9)],codeword_buf12[n*6+(16*C+9)],codeword_buf11[n*6+(16*C+9)],codeword_buf10[n*6+(16*C+9)],codeword_buf9[n*6+(16*C+9)],codeword_buf8[n*6+(16*C+9)],codeword_buf7[n*6+(16*C+9)],codeword_buf6[n*6+(16*C+9)],codeword_buf5[n*6+(16*C+9)],codeword_buf4[n*6+(16*C+9)],codeword_buf3[n*6+(16*C+9)],codeword_buf2[n*6+(16*C+9)],codeword_buf1[n*6+(16*C+9)],codeword_buf16[n*7+(16*C+9)],codeword_buf15[n*7+(16*C+9)],codeword_buf14[n*7+(16*C+9)],codeword_buf13[n*7+(16*C+9)],codeword_buf12[n*7+(16*C+9)],codeword_buf11[n*7+(16*C+9)],codeword_buf10[n*7+(16*C+9)],codeword_buf9[n*7+(16*C+9)],codeword_buf8[n*7+(16*C+9)],codeword_buf7[n*7+(16*C+9)],codeword_buf6[n*7+(16*C+9)],codeword_buf5[n*7+(16*C+9)],codeword_buf4[n*7+(16*C+9)],codeword_buf3[n*7+(16*C+9)],codeword_buf2[n*7+(16*C+9)],codeword_buf1[n*7+(16*C+9)],codeword_buf16[n*8+(16*C+9)],codeword_buf15[n*8+(16*C+9)],codeword_buf14[n*8+(16*C+9)],codeword_buf13[n*8+(16*C+9)],codeword_buf12[n*8+(16*C+9)],codeword_buf11[n*8+(16*C+9)],codeword_buf10[n*8+(16*C+9)],codeword_buf9[n*8+(16*C+9)],codeword_buf8[n*8+(16*C+9)],codeword_buf7[n*8+(16*C+9)],codeword_buf6[n*8+(16*C+9)],codeword_buf5[n*8+(16*C+9)],codeword_buf4[n*8+(16*C+9)],codeword_buf3[n*8+(16*C+9)],codeword_buf2[n*8+(16*C+9)],codeword_buf1[n*8+(16*C+9)],codeword_buf16[n*9+(16*C+9)],codeword_buf15[n*9+(16*C+9)],codeword_buf14[n*9+(16*C+9)],codeword_buf13[n*9+(16*C+9)],codeword_buf12[n*9+(16*C+9)],codeword_buf11[n*9+(16*C+9)],codeword_buf10[n*9+(16*C+9)],codeword_buf9[n*9+(16*C+9)],codeword_buf8[n*9+(16*C+9)],codeword_buf7[n*9+(16*C+9)],codeword_buf6[n*9+(16*C+9)],codeword_buf5[n*9+(16*C+9)],codeword_buf4[n*9+(16*C+9)],codeword_buf3[n*9+(16*C+9)],codeword_buf2[n*9+(16*C+9)],codeword_buf1[n*9+(16*C+9)],codeword_buf16[n*10+(16*C+9)],codeword_buf15[n*10+(16*C+9)],codeword_buf14[n*10+(16*C+9)],codeword_buf13[n*10+(16*C+9)],codeword_buf12[n*10+(16*C+9)],codeword_buf11[n*10+(16*C+9)],codeword_buf10[n*10+(16*C+9)],codeword_buf9[n*10+(16*C+9)],codeword_buf8[n*10+(16*C+9)],codeword_buf7[n*10+(16*C+9)],codeword_buf6[n*10+(16*C+9)],codeword_buf5[n*10+(16*C+9)],codeword_buf4[n*10+(16*C+9)],codeword_buf3[n*10+(16*C+9)],codeword_buf2[n*10+(16*C+9)],codeword_buf1[n*10+(16*C+9)],codeword_buf16[n*11+(16*C+9)],codeword_buf15[n*11+(16*C+9)],codeword_buf14[n*11+(16*C+9)],codeword_buf13[n*11+(16*C+9)],codeword_buf12[n*11+(16*C+9)],codeword_buf11[n*11+(16*C+9)],codeword_buf10[n*11+(16*C+9)],codeword_buf9[n*11+(16*C+9)],codeword_buf8[n*11+(16*C+9)],codeword_buf7[n*11+(16*C+9)],codeword_buf6[n*11+(16*C+9)],codeword_buf5[n*11+(16*C+9)],codeword_buf4[n*11+(16*C+9)],codeword_buf3[n*11+(16*C+9)],codeword_buf2[n*11+(16*C+9)],codeword_buf1[n*11+(16*C+9)],codeword_buf16[n*12+(16*C+9)],codeword_buf15[n*12+(16*C+9)],codeword_buf14[n*12+(16*C+9)],codeword_buf13[n*12+(16*C+9)],codeword_buf12[n*12+(16*C+9)],codeword_buf11[n*12+(16*C+9)],codeword_buf10[n*12+(16*C+9)],codeword_buf9[n*12+(16*C+9)],codeword_buf8[n*12+(16*C+9)],codeword_buf7[n*12+(16*C+9)],codeword_buf6[n*12+(16*C+9)],codeword_buf5[n*12+(16*C+9)],codeword_buf4[n*12+(16*C+9)],codeword_buf3[n*12+(16*C+9)],codeword_buf2[n*12+(16*C+9)],codeword_buf1[n*12+(16*C+9)],codeword_buf16[n*13+(16*C+9)],codeword_buf15[n*13+(16*C+9)],codeword_buf14[n*13+(16*C+9)],codeword_buf13[n*13+(16*C+9)],codeword_buf12[n*13+(16*C+9)],codeword_buf11[n*13+(16*C+9)],codeword_buf10[n*13+(16*C+9)],codeword_buf9[n*13+(16*C+9)],codeword_buf8[n*13+(16*C+9)],codeword_buf7[n*13+(16*C+9)],codeword_buf6[n*13+(16*C+9)],codeword_buf5[n*13+(16*C+9)],codeword_buf4[n*13+(16*C+9)],codeword_buf3[n*13+(16*C+9)],codeword_buf2[n*13+(16*C+9)],codeword_buf1[n*13+(16*C+9)],codeword_buf16[n*14+(16*C+9)],codeword_buf15[n*14+(16*C+9)],codeword_buf14[n*14+(16*C+9)],codeword_buf13[n*14+(16*C+9)],codeword_buf12[n*14+(16*C+9)],codeword_buf11[n*14+(16*C+9)],codeword_buf10[n*14+(16*C+9)],codeword_buf9[n*14+(16*C+9)],codeword_buf8[n*14+(16*C+9)],codeword_buf7[n*14+(16*C+9)],codeword_buf6[n*14+(16*C+9)],codeword_buf5[n*14+(16*C+9)],codeword_buf4[n*14+(16*C+9)],codeword_buf3[n*14+(16*C+9)],codeword_buf2[n*14+(16*C+9)],codeword_buf1[n*14+(16*C+9)],codeword_buf16[n*15+(16*C+9)],codeword_buf15[n*15+(16*C+9)],codeword_buf14[n*15+(16*C+9)],codeword_buf13[n*15+(16*C+9)],codeword_buf12[n*15+(16*C+9)],codeword_buf11[n*15+(16*C+9)],codeword_buf10[n*15+(16*C+9)],codeword_buf9[n*15+(16*C+9)],codeword_buf8[n*15+(16*C+9)],codeword_buf7[n*15+(16*C+9)],codeword_buf6[n*15+(16*C+9)],codeword_buf5[n*15+(16*C+9)],codeword_buf4[n*15+(16*C+9)],codeword_buf3[n*15+(16*C+9)],codeword_buf2[n*15+(16*C+9)],codeword_buf1[n*15+(16*C+9)]};
                            in_rec11 <= {codeword_buf16[n*0+(16*C+10)],codeword_buf15[n*0+(16*C+10)],codeword_buf14[n*0+(16*C+10)],codeword_buf13[n*0+(16*C+10)],codeword_buf12[n*0+(16*C+10)],codeword_buf11[n*0+(16*C+10)],codeword_buf10[n*0+(16*C+10)],codeword_buf9[n*0+(16*C+10)],codeword_buf8[n*0+(16*C+10)],codeword_buf7[n*0+(16*C+10)],codeword_buf6[n*0+(16*C+10)],codeword_buf5[n*0+(16*C+10)],codeword_buf4[n*0+(16*C+10)],codeword_buf3[n*0+(16*C+10)],codeword_buf2[n*0+(16*C+10)],codeword_buf1[n*0+(16*C+10)],codeword_buf16[n*1+(16*C+10)],codeword_buf15[n*1+(16*C+10)],codeword_buf14[n*1+(16*C+10)],codeword_buf13[n*1+(16*C+10)],codeword_buf12[n*1+(16*C+10)],codeword_buf11[n*1+(16*C+10)],codeword_buf10[n*1+(16*C+10)],codeword_buf9[n*1+(16*C+10)],codeword_buf8[n*1+(16*C+10)],codeword_buf7[n*1+(16*C+10)],codeword_buf6[n*1+(16*C+10)],codeword_buf5[n*1+(16*C+10)],codeword_buf4[n*1+(16*C+10)],codeword_buf3[n*1+(16*C+10)],codeword_buf2[n*1+(16*C+10)],codeword_buf1[n*1+(16*C+10)],codeword_buf16[n*2+(16*C+10)],codeword_buf15[n*2+(16*C+10)],codeword_buf14[n*2+(16*C+10)],codeword_buf13[n*2+(16*C+10)],codeword_buf12[n*2+(16*C+10)],codeword_buf11[n*2+(16*C+10)],codeword_buf10[n*2+(16*C+10)],codeword_buf9[n*2+(16*C+10)],codeword_buf8[n*2+(16*C+10)],codeword_buf7[n*2+(16*C+10)],codeword_buf6[n*2+(16*C+10)],codeword_buf5[n*2+(16*C+10)],codeword_buf4[n*2+(16*C+10)],codeword_buf3[n*2+(16*C+10)],codeword_buf2[n*2+(16*C+10)],codeword_buf1[n*2+(16*C+10)],codeword_buf16[n*3+(16*C+10)],codeword_buf15[n*3+(16*C+10)],codeword_buf14[n*3+(16*C+10)],codeword_buf13[n*3+(16*C+10)],codeword_buf12[n*3+(16*C+10)],codeword_buf11[n*3+(16*C+10)],codeword_buf10[n*3+(16*C+10)],codeword_buf9[n*3+(16*C+10)],codeword_buf8[n*3+(16*C+10)],codeword_buf7[n*3+(16*C+10)],codeword_buf6[n*3+(16*C+10)],codeword_buf5[n*3+(16*C+10)],codeword_buf4[n*3+(16*C+10)],codeword_buf3[n*3+(16*C+10)],codeword_buf2[n*3+(16*C+10)],codeword_buf1[n*3+(16*C+10)],codeword_buf16[n*4+(16*C+10)],codeword_buf15[n*4+(16*C+10)],codeword_buf14[n*4+(16*C+10)],codeword_buf13[n*4+(16*C+10)],codeword_buf12[n*4+(16*C+10)],codeword_buf11[n*4+(16*C+10)],codeword_buf10[n*4+(16*C+10)],codeword_buf9[n*4+(16*C+10)],codeword_buf8[n*4+(16*C+10)],codeword_buf7[n*4+(16*C+10)],codeword_buf6[n*4+(16*C+10)],codeword_buf5[n*4+(16*C+10)],codeword_buf4[n*4+(16*C+10)],codeword_buf3[n*4+(16*C+10)],codeword_buf2[n*4+(16*C+10)],codeword_buf1[n*4+(16*C+10)],codeword_buf16[n*5+(16*C+10)],codeword_buf15[n*5+(16*C+10)],codeword_buf14[n*5+(16*C+10)],codeword_buf13[n*5+(16*C+10)],codeword_buf12[n*5+(16*C+10)],codeword_buf11[n*5+(16*C+10)],codeword_buf10[n*5+(16*C+10)],codeword_buf9[n*5+(16*C+10)],codeword_buf8[n*5+(16*C+10)],codeword_buf7[n*5+(16*C+10)],codeword_buf6[n*5+(16*C+10)],codeword_buf5[n*5+(16*C+10)],codeword_buf4[n*5+(16*C+10)],codeword_buf3[n*5+(16*C+10)],codeword_buf2[n*5+(16*C+10)],codeword_buf1[n*5+(16*C+10)],codeword_buf16[n*6+(16*C+10)],codeword_buf15[n*6+(16*C+10)],codeword_buf14[n*6+(16*C+10)],codeword_buf13[n*6+(16*C+10)],codeword_buf12[n*6+(16*C+10)],codeword_buf11[n*6+(16*C+10)],codeword_buf10[n*6+(16*C+10)],codeword_buf9[n*6+(16*C+10)],codeword_buf8[n*6+(16*C+10)],codeword_buf7[n*6+(16*C+10)],codeword_buf6[n*6+(16*C+10)],codeword_buf5[n*6+(16*C+10)],codeword_buf4[n*6+(16*C+10)],codeword_buf3[n*6+(16*C+10)],codeword_buf2[n*6+(16*C+10)],codeword_buf1[n*6+(16*C+10)],codeword_buf16[n*7+(16*C+10)],codeword_buf15[n*7+(16*C+10)],codeword_buf14[n*7+(16*C+10)],codeword_buf13[n*7+(16*C+10)],codeword_buf12[n*7+(16*C+10)],codeword_buf11[n*7+(16*C+10)],codeword_buf10[n*7+(16*C+10)],codeword_buf9[n*7+(16*C+10)],codeword_buf8[n*7+(16*C+10)],codeword_buf7[n*7+(16*C+10)],codeword_buf6[n*7+(16*C+10)],codeword_buf5[n*7+(16*C+10)],codeword_buf4[n*7+(16*C+10)],codeword_buf3[n*7+(16*C+10)],codeword_buf2[n*7+(16*C+10)],codeword_buf1[n*7+(16*C+10)],codeword_buf16[n*8+(16*C+10)],codeword_buf15[n*8+(16*C+10)],codeword_buf14[n*8+(16*C+10)],codeword_buf13[n*8+(16*C+10)],codeword_buf12[n*8+(16*C+10)],codeword_buf11[n*8+(16*C+10)],codeword_buf10[n*8+(16*C+10)],codeword_buf9[n*8+(16*C+10)],codeword_buf8[n*8+(16*C+10)],codeword_buf7[n*8+(16*C+10)],codeword_buf6[n*8+(16*C+10)],codeword_buf5[n*8+(16*C+10)],codeword_buf4[n*8+(16*C+10)],codeword_buf3[n*8+(16*C+10)],codeword_buf2[n*8+(16*C+10)],codeword_buf1[n*8+(16*C+10)],codeword_buf16[n*9+(16*C+10)],codeword_buf15[n*9+(16*C+10)],codeword_buf14[n*9+(16*C+10)],codeword_buf13[n*9+(16*C+10)],codeword_buf12[n*9+(16*C+10)],codeword_buf11[n*9+(16*C+10)],codeword_buf10[n*9+(16*C+10)],codeword_buf9[n*9+(16*C+10)],codeword_buf8[n*9+(16*C+10)],codeword_buf7[n*9+(16*C+10)],codeword_buf6[n*9+(16*C+10)],codeword_buf5[n*9+(16*C+10)],codeword_buf4[n*9+(16*C+10)],codeword_buf3[n*9+(16*C+10)],codeword_buf2[n*9+(16*C+10)],codeword_buf1[n*9+(16*C+10)],codeword_buf16[n*10+(16*C+10)],codeword_buf15[n*10+(16*C+10)],codeword_buf14[n*10+(16*C+10)],codeword_buf13[n*10+(16*C+10)],codeword_buf12[n*10+(16*C+10)],codeword_buf11[n*10+(16*C+10)],codeword_buf10[n*10+(16*C+10)],codeword_buf9[n*10+(16*C+10)],codeword_buf8[n*10+(16*C+10)],codeword_buf7[n*10+(16*C+10)],codeword_buf6[n*10+(16*C+10)],codeword_buf5[n*10+(16*C+10)],codeword_buf4[n*10+(16*C+10)],codeword_buf3[n*10+(16*C+10)],codeword_buf2[n*10+(16*C+10)],codeword_buf1[n*10+(16*C+10)],codeword_buf16[n*11+(16*C+10)],codeword_buf15[n*11+(16*C+10)],codeword_buf14[n*11+(16*C+10)],codeword_buf13[n*11+(16*C+10)],codeword_buf12[n*11+(16*C+10)],codeword_buf11[n*11+(16*C+10)],codeword_buf10[n*11+(16*C+10)],codeword_buf9[n*11+(16*C+10)],codeword_buf8[n*11+(16*C+10)],codeword_buf7[n*11+(16*C+10)],codeword_buf6[n*11+(16*C+10)],codeword_buf5[n*11+(16*C+10)],codeword_buf4[n*11+(16*C+10)],codeword_buf3[n*11+(16*C+10)],codeword_buf2[n*11+(16*C+10)],codeword_buf1[n*11+(16*C+10)],codeword_buf16[n*12+(16*C+10)],codeword_buf15[n*12+(16*C+10)],codeword_buf14[n*12+(16*C+10)],codeword_buf13[n*12+(16*C+10)],codeword_buf12[n*12+(16*C+10)],codeword_buf11[n*12+(16*C+10)],codeword_buf10[n*12+(16*C+10)],codeword_buf9[n*12+(16*C+10)],codeword_buf8[n*12+(16*C+10)],codeword_buf7[n*12+(16*C+10)],codeword_buf6[n*12+(16*C+10)],codeword_buf5[n*12+(16*C+10)],codeword_buf4[n*12+(16*C+10)],codeword_buf3[n*12+(16*C+10)],codeword_buf2[n*12+(16*C+10)],codeword_buf1[n*12+(16*C+10)],codeword_buf16[n*13+(16*C+10)],codeword_buf15[n*13+(16*C+10)],codeword_buf14[n*13+(16*C+10)],codeword_buf13[n*13+(16*C+10)],codeword_buf12[n*13+(16*C+10)],codeword_buf11[n*13+(16*C+10)],codeword_buf10[n*13+(16*C+10)],codeword_buf9[n*13+(16*C+10)],codeword_buf8[n*13+(16*C+10)],codeword_buf7[n*13+(16*C+10)],codeword_buf6[n*13+(16*C+10)],codeword_buf5[n*13+(16*C+10)],codeword_buf4[n*13+(16*C+10)],codeword_buf3[n*13+(16*C+10)],codeword_buf2[n*13+(16*C+10)],codeword_buf1[n*13+(16*C+10)],codeword_buf16[n*14+(16*C+10)],codeword_buf15[n*14+(16*C+10)],codeword_buf14[n*14+(16*C+10)],codeword_buf13[n*14+(16*C+10)],codeword_buf12[n*14+(16*C+10)],codeword_buf11[n*14+(16*C+10)],codeword_buf10[n*14+(16*C+10)],codeword_buf9[n*14+(16*C+10)],codeword_buf8[n*14+(16*C+10)],codeword_buf7[n*14+(16*C+10)],codeword_buf6[n*14+(16*C+10)],codeword_buf5[n*14+(16*C+10)],codeword_buf4[n*14+(16*C+10)],codeword_buf3[n*14+(16*C+10)],codeword_buf2[n*14+(16*C+10)],codeword_buf1[n*14+(16*C+10)],codeword_buf16[n*15+(16*C+10)],codeword_buf15[n*15+(16*C+10)],codeword_buf14[n*15+(16*C+10)],codeword_buf13[n*15+(16*C+10)],codeword_buf12[n*15+(16*C+10)],codeword_buf11[n*15+(16*C+10)],codeword_buf10[n*15+(16*C+10)],codeword_buf9[n*15+(16*C+10)],codeword_buf8[n*15+(16*C+10)],codeword_buf7[n*15+(16*C+10)],codeword_buf6[n*15+(16*C+10)],codeword_buf5[n*15+(16*C+10)],codeword_buf4[n*15+(16*C+10)],codeword_buf3[n*15+(16*C+10)],codeword_buf2[n*15+(16*C+10)],codeword_buf1[n*15+(16*C+10)]};
                            in_rec12 <= {codeword_buf16[n*0+(16*C+11)],codeword_buf15[n*0+(16*C+11)],codeword_buf14[n*0+(16*C+11)],codeword_buf13[n*0+(16*C+11)],codeword_buf12[n*0+(16*C+11)],codeword_buf11[n*0+(16*C+11)],codeword_buf10[n*0+(16*C+11)],codeword_buf9[n*0+(16*C+11)],codeword_buf8[n*0+(16*C+11)],codeword_buf7[n*0+(16*C+11)],codeword_buf6[n*0+(16*C+11)],codeword_buf5[n*0+(16*C+11)],codeword_buf4[n*0+(16*C+11)],codeword_buf3[n*0+(16*C+11)],codeword_buf2[n*0+(16*C+11)],codeword_buf1[n*0+(16*C+11)],codeword_buf16[n*1+(16*C+11)],codeword_buf15[n*1+(16*C+11)],codeword_buf14[n*1+(16*C+11)],codeword_buf13[n*1+(16*C+11)],codeword_buf12[n*1+(16*C+11)],codeword_buf11[n*1+(16*C+11)],codeword_buf10[n*1+(16*C+11)],codeword_buf9[n*1+(16*C+11)],codeword_buf8[n*1+(16*C+11)],codeword_buf7[n*1+(16*C+11)],codeword_buf6[n*1+(16*C+11)],codeword_buf5[n*1+(16*C+11)],codeword_buf4[n*1+(16*C+11)],codeword_buf3[n*1+(16*C+11)],codeword_buf2[n*1+(16*C+11)],codeword_buf1[n*1+(16*C+11)],codeword_buf16[n*2+(16*C+11)],codeword_buf15[n*2+(16*C+11)],codeword_buf14[n*2+(16*C+11)],codeword_buf13[n*2+(16*C+11)],codeword_buf12[n*2+(16*C+11)],codeword_buf11[n*2+(16*C+11)],codeword_buf10[n*2+(16*C+11)],codeword_buf9[n*2+(16*C+11)],codeword_buf8[n*2+(16*C+11)],codeword_buf7[n*2+(16*C+11)],codeword_buf6[n*2+(16*C+11)],codeword_buf5[n*2+(16*C+11)],codeword_buf4[n*2+(16*C+11)],codeword_buf3[n*2+(16*C+11)],codeword_buf2[n*2+(16*C+11)],codeword_buf1[n*2+(16*C+11)],codeword_buf16[n*3+(16*C+11)],codeword_buf15[n*3+(16*C+11)],codeword_buf14[n*3+(16*C+11)],codeword_buf13[n*3+(16*C+11)],codeword_buf12[n*3+(16*C+11)],codeword_buf11[n*3+(16*C+11)],codeword_buf10[n*3+(16*C+11)],codeword_buf9[n*3+(16*C+11)],codeword_buf8[n*3+(16*C+11)],codeword_buf7[n*3+(16*C+11)],codeword_buf6[n*3+(16*C+11)],codeword_buf5[n*3+(16*C+11)],codeword_buf4[n*3+(16*C+11)],codeword_buf3[n*3+(16*C+11)],codeword_buf2[n*3+(16*C+11)],codeword_buf1[n*3+(16*C+11)],codeword_buf16[n*4+(16*C+11)],codeword_buf15[n*4+(16*C+11)],codeword_buf14[n*4+(16*C+11)],codeword_buf13[n*4+(16*C+11)],codeword_buf12[n*4+(16*C+11)],codeword_buf11[n*4+(16*C+11)],codeword_buf10[n*4+(16*C+11)],codeword_buf9[n*4+(16*C+11)],codeword_buf8[n*4+(16*C+11)],codeword_buf7[n*4+(16*C+11)],codeword_buf6[n*4+(16*C+11)],codeword_buf5[n*4+(16*C+11)],codeword_buf4[n*4+(16*C+11)],codeword_buf3[n*4+(16*C+11)],codeword_buf2[n*4+(16*C+11)],codeword_buf1[n*4+(16*C+11)],codeword_buf16[n*5+(16*C+11)],codeword_buf15[n*5+(16*C+11)],codeword_buf14[n*5+(16*C+11)],codeword_buf13[n*5+(16*C+11)],codeword_buf12[n*5+(16*C+11)],codeword_buf11[n*5+(16*C+11)],codeword_buf10[n*5+(16*C+11)],codeword_buf9[n*5+(16*C+11)],codeword_buf8[n*5+(16*C+11)],codeword_buf7[n*5+(16*C+11)],codeword_buf6[n*5+(16*C+11)],codeword_buf5[n*5+(16*C+11)],codeword_buf4[n*5+(16*C+11)],codeword_buf3[n*5+(16*C+11)],codeword_buf2[n*5+(16*C+11)],codeword_buf1[n*5+(16*C+11)],codeword_buf16[n*6+(16*C+11)],codeword_buf15[n*6+(16*C+11)],codeword_buf14[n*6+(16*C+11)],codeword_buf13[n*6+(16*C+11)],codeword_buf12[n*6+(16*C+11)],codeword_buf11[n*6+(16*C+11)],codeword_buf10[n*6+(16*C+11)],codeword_buf9[n*6+(16*C+11)],codeword_buf8[n*6+(16*C+11)],codeword_buf7[n*6+(16*C+11)],codeword_buf6[n*6+(16*C+11)],codeword_buf5[n*6+(16*C+11)],codeword_buf4[n*6+(16*C+11)],codeword_buf3[n*6+(16*C+11)],codeword_buf2[n*6+(16*C+11)],codeword_buf1[n*6+(16*C+11)],codeword_buf16[n*7+(16*C+11)],codeword_buf15[n*7+(16*C+11)],codeword_buf14[n*7+(16*C+11)],codeword_buf13[n*7+(16*C+11)],codeword_buf12[n*7+(16*C+11)],codeword_buf11[n*7+(16*C+11)],codeword_buf10[n*7+(16*C+11)],codeword_buf9[n*7+(16*C+11)],codeword_buf8[n*7+(16*C+11)],codeword_buf7[n*7+(16*C+11)],codeword_buf6[n*7+(16*C+11)],codeword_buf5[n*7+(16*C+11)],codeword_buf4[n*7+(16*C+11)],codeword_buf3[n*7+(16*C+11)],codeword_buf2[n*7+(16*C+11)],codeword_buf1[n*7+(16*C+11)],codeword_buf16[n*8+(16*C+11)],codeword_buf15[n*8+(16*C+11)],codeword_buf14[n*8+(16*C+11)],codeword_buf13[n*8+(16*C+11)],codeword_buf12[n*8+(16*C+11)],codeword_buf11[n*8+(16*C+11)],codeword_buf10[n*8+(16*C+11)],codeword_buf9[n*8+(16*C+11)],codeword_buf8[n*8+(16*C+11)],codeword_buf7[n*8+(16*C+11)],codeword_buf6[n*8+(16*C+11)],codeword_buf5[n*8+(16*C+11)],codeword_buf4[n*8+(16*C+11)],codeword_buf3[n*8+(16*C+11)],codeword_buf2[n*8+(16*C+11)],codeword_buf1[n*8+(16*C+11)],codeword_buf16[n*9+(16*C+11)],codeword_buf15[n*9+(16*C+11)],codeword_buf14[n*9+(16*C+11)],codeword_buf13[n*9+(16*C+11)],codeword_buf12[n*9+(16*C+11)],codeword_buf11[n*9+(16*C+11)],codeword_buf10[n*9+(16*C+11)],codeword_buf9[n*9+(16*C+11)],codeword_buf8[n*9+(16*C+11)],codeword_buf7[n*9+(16*C+11)],codeword_buf6[n*9+(16*C+11)],codeword_buf5[n*9+(16*C+11)],codeword_buf4[n*9+(16*C+11)],codeword_buf3[n*9+(16*C+11)],codeword_buf2[n*9+(16*C+11)],codeword_buf1[n*9+(16*C+11)],codeword_buf16[n*10+(16*C+11)],codeword_buf15[n*10+(16*C+11)],codeword_buf14[n*10+(16*C+11)],codeword_buf13[n*10+(16*C+11)],codeword_buf12[n*10+(16*C+11)],codeword_buf11[n*10+(16*C+11)],codeword_buf10[n*10+(16*C+11)],codeword_buf9[n*10+(16*C+11)],codeword_buf8[n*10+(16*C+11)],codeword_buf7[n*10+(16*C+11)],codeword_buf6[n*10+(16*C+11)],codeword_buf5[n*10+(16*C+11)],codeword_buf4[n*10+(16*C+11)],codeword_buf3[n*10+(16*C+11)],codeword_buf2[n*10+(16*C+11)],codeword_buf1[n*10+(16*C+11)],codeword_buf16[n*11+(16*C+11)],codeword_buf15[n*11+(16*C+11)],codeword_buf14[n*11+(16*C+11)],codeword_buf13[n*11+(16*C+11)],codeword_buf12[n*11+(16*C+11)],codeword_buf11[n*11+(16*C+11)],codeword_buf10[n*11+(16*C+11)],codeword_buf9[n*11+(16*C+11)],codeword_buf8[n*11+(16*C+11)],codeword_buf7[n*11+(16*C+11)],codeword_buf6[n*11+(16*C+11)],codeword_buf5[n*11+(16*C+11)],codeword_buf4[n*11+(16*C+11)],codeword_buf3[n*11+(16*C+11)],codeword_buf2[n*11+(16*C+11)],codeword_buf1[n*11+(16*C+11)],codeword_buf16[n*12+(16*C+11)],codeword_buf15[n*12+(16*C+11)],codeword_buf14[n*12+(16*C+11)],codeword_buf13[n*12+(16*C+11)],codeword_buf12[n*12+(16*C+11)],codeword_buf11[n*12+(16*C+11)],codeword_buf10[n*12+(16*C+11)],codeword_buf9[n*12+(16*C+11)],codeword_buf8[n*12+(16*C+11)],codeword_buf7[n*12+(16*C+11)],codeword_buf6[n*12+(16*C+11)],codeword_buf5[n*12+(16*C+11)],codeword_buf4[n*12+(16*C+11)],codeword_buf3[n*12+(16*C+11)],codeword_buf2[n*12+(16*C+11)],codeword_buf1[n*12+(16*C+11)],codeword_buf16[n*13+(16*C+11)],codeword_buf15[n*13+(16*C+11)],codeword_buf14[n*13+(16*C+11)],codeword_buf13[n*13+(16*C+11)],codeword_buf12[n*13+(16*C+11)],codeword_buf11[n*13+(16*C+11)],codeword_buf10[n*13+(16*C+11)],codeword_buf9[n*13+(16*C+11)],codeword_buf8[n*13+(16*C+11)],codeword_buf7[n*13+(16*C+11)],codeword_buf6[n*13+(16*C+11)],codeword_buf5[n*13+(16*C+11)],codeword_buf4[n*13+(16*C+11)],codeword_buf3[n*13+(16*C+11)],codeword_buf2[n*13+(16*C+11)],codeword_buf1[n*13+(16*C+11)],codeword_buf16[n*14+(16*C+11)],codeword_buf15[n*14+(16*C+11)],codeword_buf14[n*14+(16*C+11)],codeword_buf13[n*14+(16*C+11)],codeword_buf12[n*14+(16*C+11)],codeword_buf11[n*14+(16*C+11)],codeword_buf10[n*14+(16*C+11)],codeword_buf9[n*14+(16*C+11)],codeword_buf8[n*14+(16*C+11)],codeword_buf7[n*14+(16*C+11)],codeword_buf6[n*14+(16*C+11)],codeword_buf5[n*14+(16*C+11)],codeword_buf4[n*14+(16*C+11)],codeword_buf3[n*14+(16*C+11)],codeword_buf2[n*14+(16*C+11)],codeword_buf1[n*14+(16*C+11)],codeword_buf16[n*15+(16*C+11)],codeword_buf15[n*15+(16*C+11)],codeword_buf14[n*15+(16*C+11)],codeword_buf13[n*15+(16*C+11)],codeword_buf12[n*15+(16*C+11)],codeword_buf11[n*15+(16*C+11)],codeword_buf10[n*15+(16*C+11)],codeword_buf9[n*15+(16*C+11)],codeword_buf8[n*15+(16*C+11)],codeword_buf7[n*15+(16*C+11)],codeword_buf6[n*15+(16*C+11)],codeword_buf5[n*15+(16*C+11)],codeword_buf4[n*15+(16*C+11)],codeword_buf3[n*15+(16*C+11)],codeword_buf2[n*15+(16*C+11)],codeword_buf1[n*15+(16*C+11)]};
                            in_rec13 <= {codeword_buf16[n*0+(16*C+12)],codeword_buf15[n*0+(16*C+12)],codeword_buf14[n*0+(16*C+12)],codeword_buf13[n*0+(16*C+12)],codeword_buf12[n*0+(16*C+12)],codeword_buf11[n*0+(16*C+12)],codeword_buf10[n*0+(16*C+12)],codeword_buf9[n*0+(16*C+12)],codeword_buf8[n*0+(16*C+12)],codeword_buf7[n*0+(16*C+12)],codeword_buf6[n*0+(16*C+12)],codeword_buf5[n*0+(16*C+12)],codeword_buf4[n*0+(16*C+12)],codeword_buf3[n*0+(16*C+12)],codeword_buf2[n*0+(16*C+12)],codeword_buf1[n*0+(16*C+12)],codeword_buf16[n*1+(16*C+12)],codeword_buf15[n*1+(16*C+12)],codeword_buf14[n*1+(16*C+12)],codeword_buf13[n*1+(16*C+12)],codeword_buf12[n*1+(16*C+12)],codeword_buf11[n*1+(16*C+12)],codeword_buf10[n*1+(16*C+12)],codeword_buf9[n*1+(16*C+12)],codeword_buf8[n*1+(16*C+12)],codeword_buf7[n*1+(16*C+12)],codeword_buf6[n*1+(16*C+12)],codeword_buf5[n*1+(16*C+12)],codeword_buf4[n*1+(16*C+12)],codeword_buf3[n*1+(16*C+12)],codeword_buf2[n*1+(16*C+12)],codeword_buf1[n*1+(16*C+12)],codeword_buf16[n*2+(16*C+12)],codeword_buf15[n*2+(16*C+12)],codeword_buf14[n*2+(16*C+12)],codeword_buf13[n*2+(16*C+12)],codeword_buf12[n*2+(16*C+12)],codeword_buf11[n*2+(16*C+12)],codeword_buf10[n*2+(16*C+12)],codeword_buf9[n*2+(16*C+12)],codeword_buf8[n*2+(16*C+12)],codeword_buf7[n*2+(16*C+12)],codeword_buf6[n*2+(16*C+12)],codeword_buf5[n*2+(16*C+12)],codeword_buf4[n*2+(16*C+12)],codeword_buf3[n*2+(16*C+12)],codeword_buf2[n*2+(16*C+12)],codeword_buf1[n*2+(16*C+12)],codeword_buf16[n*3+(16*C+12)],codeword_buf15[n*3+(16*C+12)],codeword_buf14[n*3+(16*C+12)],codeword_buf13[n*3+(16*C+12)],codeword_buf12[n*3+(16*C+12)],codeword_buf11[n*3+(16*C+12)],codeword_buf10[n*3+(16*C+12)],codeword_buf9[n*3+(16*C+12)],codeword_buf8[n*3+(16*C+12)],codeword_buf7[n*3+(16*C+12)],codeword_buf6[n*3+(16*C+12)],codeword_buf5[n*3+(16*C+12)],codeword_buf4[n*3+(16*C+12)],codeword_buf3[n*3+(16*C+12)],codeword_buf2[n*3+(16*C+12)],codeword_buf1[n*3+(16*C+12)],codeword_buf16[n*4+(16*C+12)],codeword_buf15[n*4+(16*C+12)],codeword_buf14[n*4+(16*C+12)],codeword_buf13[n*4+(16*C+12)],codeword_buf12[n*4+(16*C+12)],codeword_buf11[n*4+(16*C+12)],codeword_buf10[n*4+(16*C+12)],codeword_buf9[n*4+(16*C+12)],codeword_buf8[n*4+(16*C+12)],codeword_buf7[n*4+(16*C+12)],codeword_buf6[n*4+(16*C+12)],codeword_buf5[n*4+(16*C+12)],codeword_buf4[n*4+(16*C+12)],codeword_buf3[n*4+(16*C+12)],codeword_buf2[n*4+(16*C+12)],codeword_buf1[n*4+(16*C+12)],codeword_buf16[n*5+(16*C+12)],codeword_buf15[n*5+(16*C+12)],codeword_buf14[n*5+(16*C+12)],codeword_buf13[n*5+(16*C+12)],codeword_buf12[n*5+(16*C+12)],codeword_buf11[n*5+(16*C+12)],codeword_buf10[n*5+(16*C+12)],codeword_buf9[n*5+(16*C+12)],codeword_buf8[n*5+(16*C+12)],codeword_buf7[n*5+(16*C+12)],codeword_buf6[n*5+(16*C+12)],codeword_buf5[n*5+(16*C+12)],codeword_buf4[n*5+(16*C+12)],codeword_buf3[n*5+(16*C+12)],codeword_buf2[n*5+(16*C+12)],codeword_buf1[n*5+(16*C+12)],codeword_buf16[n*6+(16*C+12)],codeword_buf15[n*6+(16*C+12)],codeword_buf14[n*6+(16*C+12)],codeword_buf13[n*6+(16*C+12)],codeword_buf12[n*6+(16*C+12)],codeword_buf11[n*6+(16*C+12)],codeword_buf10[n*6+(16*C+12)],codeword_buf9[n*6+(16*C+12)],codeword_buf8[n*6+(16*C+12)],codeword_buf7[n*6+(16*C+12)],codeword_buf6[n*6+(16*C+12)],codeword_buf5[n*6+(16*C+12)],codeword_buf4[n*6+(16*C+12)],codeword_buf3[n*6+(16*C+12)],codeword_buf2[n*6+(16*C+12)],codeword_buf1[n*6+(16*C+12)],codeword_buf16[n*7+(16*C+12)],codeword_buf15[n*7+(16*C+12)],codeword_buf14[n*7+(16*C+12)],codeword_buf13[n*7+(16*C+12)],codeword_buf12[n*7+(16*C+12)],codeword_buf11[n*7+(16*C+12)],codeword_buf10[n*7+(16*C+12)],codeword_buf9[n*7+(16*C+12)],codeword_buf8[n*7+(16*C+12)],codeword_buf7[n*7+(16*C+12)],codeword_buf6[n*7+(16*C+12)],codeword_buf5[n*7+(16*C+12)],codeword_buf4[n*7+(16*C+12)],codeword_buf3[n*7+(16*C+12)],codeword_buf2[n*7+(16*C+12)],codeword_buf1[n*7+(16*C+12)],codeword_buf16[n*8+(16*C+12)],codeword_buf15[n*8+(16*C+12)],codeword_buf14[n*8+(16*C+12)],codeword_buf13[n*8+(16*C+12)],codeword_buf12[n*8+(16*C+12)],codeword_buf11[n*8+(16*C+12)],codeword_buf10[n*8+(16*C+12)],codeword_buf9[n*8+(16*C+12)],codeword_buf8[n*8+(16*C+12)],codeword_buf7[n*8+(16*C+12)],codeword_buf6[n*8+(16*C+12)],codeword_buf5[n*8+(16*C+12)],codeword_buf4[n*8+(16*C+12)],codeword_buf3[n*8+(16*C+12)],codeword_buf2[n*8+(16*C+12)],codeword_buf1[n*8+(16*C+12)],codeword_buf16[n*9+(16*C+12)],codeword_buf15[n*9+(16*C+12)],codeword_buf14[n*9+(16*C+12)],codeword_buf13[n*9+(16*C+12)],codeword_buf12[n*9+(16*C+12)],codeword_buf11[n*9+(16*C+12)],codeword_buf10[n*9+(16*C+12)],codeword_buf9[n*9+(16*C+12)],codeword_buf8[n*9+(16*C+12)],codeword_buf7[n*9+(16*C+12)],codeword_buf6[n*9+(16*C+12)],codeword_buf5[n*9+(16*C+12)],codeword_buf4[n*9+(16*C+12)],codeword_buf3[n*9+(16*C+12)],codeword_buf2[n*9+(16*C+12)],codeword_buf1[n*9+(16*C+12)],codeword_buf16[n*10+(16*C+12)],codeword_buf15[n*10+(16*C+12)],codeword_buf14[n*10+(16*C+12)],codeword_buf13[n*10+(16*C+12)],codeword_buf12[n*10+(16*C+12)],codeword_buf11[n*10+(16*C+12)],codeword_buf10[n*10+(16*C+12)],codeword_buf9[n*10+(16*C+12)],codeword_buf8[n*10+(16*C+12)],codeword_buf7[n*10+(16*C+12)],codeword_buf6[n*10+(16*C+12)],codeword_buf5[n*10+(16*C+12)],codeword_buf4[n*10+(16*C+12)],codeword_buf3[n*10+(16*C+12)],codeword_buf2[n*10+(16*C+12)],codeword_buf1[n*10+(16*C+12)],codeword_buf16[n*11+(16*C+12)],codeword_buf15[n*11+(16*C+12)],codeword_buf14[n*11+(16*C+12)],codeword_buf13[n*11+(16*C+12)],codeword_buf12[n*11+(16*C+12)],codeword_buf11[n*11+(16*C+12)],codeword_buf10[n*11+(16*C+12)],codeword_buf9[n*11+(16*C+12)],codeword_buf8[n*11+(16*C+12)],codeword_buf7[n*11+(16*C+12)],codeword_buf6[n*11+(16*C+12)],codeword_buf5[n*11+(16*C+12)],codeword_buf4[n*11+(16*C+12)],codeword_buf3[n*11+(16*C+12)],codeword_buf2[n*11+(16*C+12)],codeword_buf1[n*11+(16*C+12)],codeword_buf16[n*12+(16*C+12)],codeword_buf15[n*12+(16*C+12)],codeword_buf14[n*12+(16*C+12)],codeword_buf13[n*12+(16*C+12)],codeword_buf12[n*12+(16*C+12)],codeword_buf11[n*12+(16*C+12)],codeword_buf10[n*12+(16*C+12)],codeword_buf9[n*12+(16*C+12)],codeword_buf8[n*12+(16*C+12)],codeword_buf7[n*12+(16*C+12)],codeword_buf6[n*12+(16*C+12)],codeword_buf5[n*12+(16*C+12)],codeword_buf4[n*12+(16*C+12)],codeword_buf3[n*12+(16*C+12)],codeword_buf2[n*12+(16*C+12)],codeword_buf1[n*12+(16*C+12)],codeword_buf16[n*13+(16*C+12)],codeword_buf15[n*13+(16*C+12)],codeword_buf14[n*13+(16*C+12)],codeword_buf13[n*13+(16*C+12)],codeword_buf12[n*13+(16*C+12)],codeword_buf11[n*13+(16*C+12)],codeword_buf10[n*13+(16*C+12)],codeword_buf9[n*13+(16*C+12)],codeword_buf8[n*13+(16*C+12)],codeword_buf7[n*13+(16*C+12)],codeword_buf6[n*13+(16*C+12)],codeword_buf5[n*13+(16*C+12)],codeword_buf4[n*13+(16*C+12)],codeword_buf3[n*13+(16*C+12)],codeword_buf2[n*13+(16*C+12)],codeword_buf1[n*13+(16*C+12)],codeword_buf16[n*14+(16*C+12)],codeword_buf15[n*14+(16*C+12)],codeword_buf14[n*14+(16*C+12)],codeword_buf13[n*14+(16*C+12)],codeword_buf12[n*14+(16*C+12)],codeword_buf11[n*14+(16*C+12)],codeword_buf10[n*14+(16*C+12)],codeword_buf9[n*14+(16*C+12)],codeword_buf8[n*14+(16*C+12)],codeword_buf7[n*14+(16*C+12)],codeword_buf6[n*14+(16*C+12)],codeword_buf5[n*14+(16*C+12)],codeword_buf4[n*14+(16*C+12)],codeword_buf3[n*14+(16*C+12)],codeword_buf2[n*14+(16*C+12)],codeword_buf1[n*14+(16*C+12)],codeword_buf16[n*15+(16*C+12)],codeword_buf15[n*15+(16*C+12)],codeword_buf14[n*15+(16*C+12)],codeword_buf13[n*15+(16*C+12)],codeword_buf12[n*15+(16*C+12)],codeword_buf11[n*15+(16*C+12)],codeword_buf10[n*15+(16*C+12)],codeword_buf9[n*15+(16*C+12)],codeword_buf8[n*15+(16*C+12)],codeword_buf7[n*15+(16*C+12)],codeword_buf6[n*15+(16*C+12)],codeword_buf5[n*15+(16*C+12)],codeword_buf4[n*15+(16*C+12)],codeword_buf3[n*15+(16*C+12)],codeword_buf2[n*15+(16*C+12)],codeword_buf1[n*15+(16*C+12)]};
                            in_rec14 <= {codeword_buf16[n*0+(16*C+13)],codeword_buf15[n*0+(16*C+13)],codeword_buf14[n*0+(16*C+13)],codeword_buf13[n*0+(16*C+13)],codeword_buf12[n*0+(16*C+13)],codeword_buf11[n*0+(16*C+13)],codeword_buf10[n*0+(16*C+13)],codeword_buf9[n*0+(16*C+13)],codeword_buf8[n*0+(16*C+13)],codeword_buf7[n*0+(16*C+13)],codeword_buf6[n*0+(16*C+13)],codeword_buf5[n*0+(16*C+13)],codeword_buf4[n*0+(16*C+13)],codeword_buf3[n*0+(16*C+13)],codeword_buf2[n*0+(16*C+13)],codeword_buf1[n*0+(16*C+13)],codeword_buf16[n*1+(16*C+13)],codeword_buf15[n*1+(16*C+13)],codeword_buf14[n*1+(16*C+13)],codeword_buf13[n*1+(16*C+13)],codeword_buf12[n*1+(16*C+13)],codeword_buf11[n*1+(16*C+13)],codeword_buf10[n*1+(16*C+13)],codeword_buf9[n*1+(16*C+13)],codeword_buf8[n*1+(16*C+13)],codeword_buf7[n*1+(16*C+13)],codeword_buf6[n*1+(16*C+13)],codeword_buf5[n*1+(16*C+13)],codeword_buf4[n*1+(16*C+13)],codeword_buf3[n*1+(16*C+13)],codeword_buf2[n*1+(16*C+13)],codeword_buf1[n*1+(16*C+13)],codeword_buf16[n*2+(16*C+13)],codeword_buf15[n*2+(16*C+13)],codeword_buf14[n*2+(16*C+13)],codeword_buf13[n*2+(16*C+13)],codeword_buf12[n*2+(16*C+13)],codeword_buf11[n*2+(16*C+13)],codeword_buf10[n*2+(16*C+13)],codeword_buf9[n*2+(16*C+13)],codeword_buf8[n*2+(16*C+13)],codeword_buf7[n*2+(16*C+13)],codeword_buf6[n*2+(16*C+13)],codeword_buf5[n*2+(16*C+13)],codeword_buf4[n*2+(16*C+13)],codeword_buf3[n*2+(16*C+13)],codeword_buf2[n*2+(16*C+13)],codeword_buf1[n*2+(16*C+13)],codeword_buf16[n*3+(16*C+13)],codeword_buf15[n*3+(16*C+13)],codeword_buf14[n*3+(16*C+13)],codeword_buf13[n*3+(16*C+13)],codeword_buf12[n*3+(16*C+13)],codeword_buf11[n*3+(16*C+13)],codeword_buf10[n*3+(16*C+13)],codeword_buf9[n*3+(16*C+13)],codeword_buf8[n*3+(16*C+13)],codeword_buf7[n*3+(16*C+13)],codeword_buf6[n*3+(16*C+13)],codeword_buf5[n*3+(16*C+13)],codeword_buf4[n*3+(16*C+13)],codeword_buf3[n*3+(16*C+13)],codeword_buf2[n*3+(16*C+13)],codeword_buf1[n*3+(16*C+13)],codeword_buf16[n*4+(16*C+13)],codeword_buf15[n*4+(16*C+13)],codeword_buf14[n*4+(16*C+13)],codeword_buf13[n*4+(16*C+13)],codeword_buf12[n*4+(16*C+13)],codeword_buf11[n*4+(16*C+13)],codeword_buf10[n*4+(16*C+13)],codeword_buf9[n*4+(16*C+13)],codeword_buf8[n*4+(16*C+13)],codeword_buf7[n*4+(16*C+13)],codeword_buf6[n*4+(16*C+13)],codeword_buf5[n*4+(16*C+13)],codeword_buf4[n*4+(16*C+13)],codeword_buf3[n*4+(16*C+13)],codeword_buf2[n*4+(16*C+13)],codeword_buf1[n*4+(16*C+13)],codeword_buf16[n*5+(16*C+13)],codeword_buf15[n*5+(16*C+13)],codeword_buf14[n*5+(16*C+13)],codeword_buf13[n*5+(16*C+13)],codeword_buf12[n*5+(16*C+13)],codeword_buf11[n*5+(16*C+13)],codeword_buf10[n*5+(16*C+13)],codeword_buf9[n*5+(16*C+13)],codeword_buf8[n*5+(16*C+13)],codeword_buf7[n*5+(16*C+13)],codeword_buf6[n*5+(16*C+13)],codeword_buf5[n*5+(16*C+13)],codeword_buf4[n*5+(16*C+13)],codeword_buf3[n*5+(16*C+13)],codeword_buf2[n*5+(16*C+13)],codeword_buf1[n*5+(16*C+13)],codeword_buf16[n*6+(16*C+13)],codeword_buf15[n*6+(16*C+13)],codeword_buf14[n*6+(16*C+13)],codeword_buf13[n*6+(16*C+13)],codeword_buf12[n*6+(16*C+13)],codeword_buf11[n*6+(16*C+13)],codeword_buf10[n*6+(16*C+13)],codeword_buf9[n*6+(16*C+13)],codeword_buf8[n*6+(16*C+13)],codeword_buf7[n*6+(16*C+13)],codeword_buf6[n*6+(16*C+13)],codeword_buf5[n*6+(16*C+13)],codeword_buf4[n*6+(16*C+13)],codeword_buf3[n*6+(16*C+13)],codeword_buf2[n*6+(16*C+13)],codeword_buf1[n*6+(16*C+13)],codeword_buf16[n*7+(16*C+13)],codeword_buf15[n*7+(16*C+13)],codeword_buf14[n*7+(16*C+13)],codeword_buf13[n*7+(16*C+13)],codeword_buf12[n*7+(16*C+13)],codeword_buf11[n*7+(16*C+13)],codeword_buf10[n*7+(16*C+13)],codeword_buf9[n*7+(16*C+13)],codeword_buf8[n*7+(16*C+13)],codeword_buf7[n*7+(16*C+13)],codeword_buf6[n*7+(16*C+13)],codeword_buf5[n*7+(16*C+13)],codeword_buf4[n*7+(16*C+13)],codeword_buf3[n*7+(16*C+13)],codeword_buf2[n*7+(16*C+13)],codeword_buf1[n*7+(16*C+13)],codeword_buf16[n*8+(16*C+13)],codeword_buf15[n*8+(16*C+13)],codeword_buf14[n*8+(16*C+13)],codeword_buf13[n*8+(16*C+13)],codeword_buf12[n*8+(16*C+13)],codeword_buf11[n*8+(16*C+13)],codeword_buf10[n*8+(16*C+13)],codeword_buf9[n*8+(16*C+13)],codeword_buf8[n*8+(16*C+13)],codeword_buf7[n*8+(16*C+13)],codeword_buf6[n*8+(16*C+13)],codeword_buf5[n*8+(16*C+13)],codeword_buf4[n*8+(16*C+13)],codeword_buf3[n*8+(16*C+13)],codeword_buf2[n*8+(16*C+13)],codeword_buf1[n*8+(16*C+13)],codeword_buf16[n*9+(16*C+13)],codeword_buf15[n*9+(16*C+13)],codeword_buf14[n*9+(16*C+13)],codeword_buf13[n*9+(16*C+13)],codeword_buf12[n*9+(16*C+13)],codeword_buf11[n*9+(16*C+13)],codeword_buf10[n*9+(16*C+13)],codeword_buf9[n*9+(16*C+13)],codeword_buf8[n*9+(16*C+13)],codeword_buf7[n*9+(16*C+13)],codeword_buf6[n*9+(16*C+13)],codeword_buf5[n*9+(16*C+13)],codeword_buf4[n*9+(16*C+13)],codeword_buf3[n*9+(16*C+13)],codeword_buf2[n*9+(16*C+13)],codeword_buf1[n*9+(16*C+13)],codeword_buf16[n*10+(16*C+13)],codeword_buf15[n*10+(16*C+13)],codeword_buf14[n*10+(16*C+13)],codeword_buf13[n*10+(16*C+13)],codeword_buf12[n*10+(16*C+13)],codeword_buf11[n*10+(16*C+13)],codeword_buf10[n*10+(16*C+13)],codeword_buf9[n*10+(16*C+13)],codeword_buf8[n*10+(16*C+13)],codeword_buf7[n*10+(16*C+13)],codeword_buf6[n*10+(16*C+13)],codeword_buf5[n*10+(16*C+13)],codeword_buf4[n*10+(16*C+13)],codeword_buf3[n*10+(16*C+13)],codeword_buf2[n*10+(16*C+13)],codeword_buf1[n*10+(16*C+13)],codeword_buf16[n*11+(16*C+13)],codeword_buf15[n*11+(16*C+13)],codeword_buf14[n*11+(16*C+13)],codeword_buf13[n*11+(16*C+13)],codeword_buf12[n*11+(16*C+13)],codeword_buf11[n*11+(16*C+13)],codeword_buf10[n*11+(16*C+13)],codeword_buf9[n*11+(16*C+13)],codeword_buf8[n*11+(16*C+13)],codeword_buf7[n*11+(16*C+13)],codeword_buf6[n*11+(16*C+13)],codeword_buf5[n*11+(16*C+13)],codeword_buf4[n*11+(16*C+13)],codeword_buf3[n*11+(16*C+13)],codeword_buf2[n*11+(16*C+13)],codeword_buf1[n*11+(16*C+13)],codeword_buf16[n*12+(16*C+13)],codeword_buf15[n*12+(16*C+13)],codeword_buf14[n*12+(16*C+13)],codeword_buf13[n*12+(16*C+13)],codeword_buf12[n*12+(16*C+13)],codeword_buf11[n*12+(16*C+13)],codeword_buf10[n*12+(16*C+13)],codeword_buf9[n*12+(16*C+13)],codeword_buf8[n*12+(16*C+13)],codeword_buf7[n*12+(16*C+13)],codeword_buf6[n*12+(16*C+13)],codeword_buf5[n*12+(16*C+13)],codeword_buf4[n*12+(16*C+13)],codeword_buf3[n*12+(16*C+13)],codeword_buf2[n*12+(16*C+13)],codeword_buf1[n*12+(16*C+13)],codeword_buf16[n*13+(16*C+13)],codeword_buf15[n*13+(16*C+13)],codeword_buf14[n*13+(16*C+13)],codeword_buf13[n*13+(16*C+13)],codeword_buf12[n*13+(16*C+13)],codeword_buf11[n*13+(16*C+13)],codeword_buf10[n*13+(16*C+13)],codeword_buf9[n*13+(16*C+13)],codeword_buf8[n*13+(16*C+13)],codeword_buf7[n*13+(16*C+13)],codeword_buf6[n*13+(16*C+13)],codeword_buf5[n*13+(16*C+13)],codeword_buf4[n*13+(16*C+13)],codeword_buf3[n*13+(16*C+13)],codeword_buf2[n*13+(16*C+13)],codeword_buf1[n*13+(16*C+13)],codeword_buf16[n*14+(16*C+13)],codeword_buf15[n*14+(16*C+13)],codeword_buf14[n*14+(16*C+13)],codeword_buf13[n*14+(16*C+13)],codeword_buf12[n*14+(16*C+13)],codeword_buf11[n*14+(16*C+13)],codeword_buf10[n*14+(16*C+13)],codeword_buf9[n*14+(16*C+13)],codeword_buf8[n*14+(16*C+13)],codeword_buf7[n*14+(16*C+13)],codeword_buf6[n*14+(16*C+13)],codeword_buf5[n*14+(16*C+13)],codeword_buf4[n*14+(16*C+13)],codeword_buf3[n*14+(16*C+13)],codeword_buf2[n*14+(16*C+13)],codeword_buf1[n*14+(16*C+13)],codeword_buf16[n*15+(16*C+13)],codeword_buf15[n*15+(16*C+13)],codeword_buf14[n*15+(16*C+13)],codeword_buf13[n*15+(16*C+13)],codeword_buf12[n*15+(16*C+13)],codeword_buf11[n*15+(16*C+13)],codeword_buf10[n*15+(16*C+13)],codeword_buf9[n*15+(16*C+13)],codeword_buf8[n*15+(16*C+13)],codeword_buf7[n*15+(16*C+13)],codeword_buf6[n*15+(16*C+13)],codeword_buf5[n*15+(16*C+13)],codeword_buf4[n*15+(16*C+13)],codeword_buf3[n*15+(16*C+13)],codeword_buf2[n*15+(16*C+13)],codeword_buf1[n*15+(16*C+13)]};
                            in_rec15 <= {codeword_buf16[n*0+(16*C+14)],codeword_buf15[n*0+(16*C+14)],codeword_buf14[n*0+(16*C+14)],codeword_buf13[n*0+(16*C+14)],codeword_buf12[n*0+(16*C+14)],codeword_buf11[n*0+(16*C+14)],codeword_buf10[n*0+(16*C+14)],codeword_buf9[n*0+(16*C+14)],codeword_buf8[n*0+(16*C+14)],codeword_buf7[n*0+(16*C+14)],codeword_buf6[n*0+(16*C+14)],codeword_buf5[n*0+(16*C+14)],codeword_buf4[n*0+(16*C+14)],codeword_buf3[n*0+(16*C+14)],codeword_buf2[n*0+(16*C+14)],codeword_buf1[n*0+(16*C+14)],codeword_buf16[n*1+(16*C+14)],codeword_buf15[n*1+(16*C+14)],codeword_buf14[n*1+(16*C+14)],codeword_buf13[n*1+(16*C+14)],codeword_buf12[n*1+(16*C+14)],codeword_buf11[n*1+(16*C+14)],codeword_buf10[n*1+(16*C+14)],codeword_buf9[n*1+(16*C+14)],codeword_buf8[n*1+(16*C+14)],codeword_buf7[n*1+(16*C+14)],codeword_buf6[n*1+(16*C+14)],codeword_buf5[n*1+(16*C+14)],codeword_buf4[n*1+(16*C+14)],codeword_buf3[n*1+(16*C+14)],codeword_buf2[n*1+(16*C+14)],codeword_buf1[n*1+(16*C+14)],codeword_buf16[n*2+(16*C+14)],codeword_buf15[n*2+(16*C+14)],codeword_buf14[n*2+(16*C+14)],codeword_buf13[n*2+(16*C+14)],codeword_buf12[n*2+(16*C+14)],codeword_buf11[n*2+(16*C+14)],codeword_buf10[n*2+(16*C+14)],codeword_buf9[n*2+(16*C+14)],codeword_buf8[n*2+(16*C+14)],codeword_buf7[n*2+(16*C+14)],codeword_buf6[n*2+(16*C+14)],codeword_buf5[n*2+(16*C+14)],codeword_buf4[n*2+(16*C+14)],codeword_buf3[n*2+(16*C+14)],codeword_buf2[n*2+(16*C+14)],codeword_buf1[n*2+(16*C+14)],codeword_buf16[n*3+(16*C+14)],codeword_buf15[n*3+(16*C+14)],codeword_buf14[n*3+(16*C+14)],codeword_buf13[n*3+(16*C+14)],codeword_buf12[n*3+(16*C+14)],codeword_buf11[n*3+(16*C+14)],codeword_buf10[n*3+(16*C+14)],codeword_buf9[n*3+(16*C+14)],codeword_buf8[n*3+(16*C+14)],codeword_buf7[n*3+(16*C+14)],codeword_buf6[n*3+(16*C+14)],codeword_buf5[n*3+(16*C+14)],codeword_buf4[n*3+(16*C+14)],codeword_buf3[n*3+(16*C+14)],codeword_buf2[n*3+(16*C+14)],codeword_buf1[n*3+(16*C+14)],codeword_buf16[n*4+(16*C+14)],codeword_buf15[n*4+(16*C+14)],codeword_buf14[n*4+(16*C+14)],codeword_buf13[n*4+(16*C+14)],codeword_buf12[n*4+(16*C+14)],codeword_buf11[n*4+(16*C+14)],codeword_buf10[n*4+(16*C+14)],codeword_buf9[n*4+(16*C+14)],codeword_buf8[n*4+(16*C+14)],codeword_buf7[n*4+(16*C+14)],codeword_buf6[n*4+(16*C+14)],codeword_buf5[n*4+(16*C+14)],codeword_buf4[n*4+(16*C+14)],codeword_buf3[n*4+(16*C+14)],codeword_buf2[n*4+(16*C+14)],codeword_buf1[n*4+(16*C+14)],codeword_buf16[n*5+(16*C+14)],codeword_buf15[n*5+(16*C+14)],codeword_buf14[n*5+(16*C+14)],codeword_buf13[n*5+(16*C+14)],codeword_buf12[n*5+(16*C+14)],codeword_buf11[n*5+(16*C+14)],codeword_buf10[n*5+(16*C+14)],codeword_buf9[n*5+(16*C+14)],codeword_buf8[n*5+(16*C+14)],codeword_buf7[n*5+(16*C+14)],codeword_buf6[n*5+(16*C+14)],codeword_buf5[n*5+(16*C+14)],codeword_buf4[n*5+(16*C+14)],codeword_buf3[n*5+(16*C+14)],codeword_buf2[n*5+(16*C+14)],codeword_buf1[n*5+(16*C+14)],codeword_buf16[n*6+(16*C+14)],codeword_buf15[n*6+(16*C+14)],codeword_buf14[n*6+(16*C+14)],codeword_buf13[n*6+(16*C+14)],codeword_buf12[n*6+(16*C+14)],codeword_buf11[n*6+(16*C+14)],codeword_buf10[n*6+(16*C+14)],codeword_buf9[n*6+(16*C+14)],codeword_buf8[n*6+(16*C+14)],codeword_buf7[n*6+(16*C+14)],codeword_buf6[n*6+(16*C+14)],codeword_buf5[n*6+(16*C+14)],codeword_buf4[n*6+(16*C+14)],codeword_buf3[n*6+(16*C+14)],codeword_buf2[n*6+(16*C+14)],codeword_buf1[n*6+(16*C+14)],codeword_buf16[n*7+(16*C+14)],codeword_buf15[n*7+(16*C+14)],codeword_buf14[n*7+(16*C+14)],codeword_buf13[n*7+(16*C+14)],codeword_buf12[n*7+(16*C+14)],codeword_buf11[n*7+(16*C+14)],codeword_buf10[n*7+(16*C+14)],codeword_buf9[n*7+(16*C+14)],codeword_buf8[n*7+(16*C+14)],codeword_buf7[n*7+(16*C+14)],codeword_buf6[n*7+(16*C+14)],codeword_buf5[n*7+(16*C+14)],codeword_buf4[n*7+(16*C+14)],codeword_buf3[n*7+(16*C+14)],codeword_buf2[n*7+(16*C+14)],codeword_buf1[n*7+(16*C+14)],codeword_buf16[n*8+(16*C+14)],codeword_buf15[n*8+(16*C+14)],codeword_buf14[n*8+(16*C+14)],codeword_buf13[n*8+(16*C+14)],codeword_buf12[n*8+(16*C+14)],codeword_buf11[n*8+(16*C+14)],codeword_buf10[n*8+(16*C+14)],codeword_buf9[n*8+(16*C+14)],codeword_buf8[n*8+(16*C+14)],codeword_buf7[n*8+(16*C+14)],codeword_buf6[n*8+(16*C+14)],codeword_buf5[n*8+(16*C+14)],codeword_buf4[n*8+(16*C+14)],codeword_buf3[n*8+(16*C+14)],codeword_buf2[n*8+(16*C+14)],codeword_buf1[n*8+(16*C+14)],codeword_buf16[n*9+(16*C+14)],codeword_buf15[n*9+(16*C+14)],codeword_buf14[n*9+(16*C+14)],codeword_buf13[n*9+(16*C+14)],codeword_buf12[n*9+(16*C+14)],codeword_buf11[n*9+(16*C+14)],codeword_buf10[n*9+(16*C+14)],codeword_buf9[n*9+(16*C+14)],codeword_buf8[n*9+(16*C+14)],codeword_buf7[n*9+(16*C+14)],codeword_buf6[n*9+(16*C+14)],codeword_buf5[n*9+(16*C+14)],codeword_buf4[n*9+(16*C+14)],codeword_buf3[n*9+(16*C+14)],codeword_buf2[n*9+(16*C+14)],codeword_buf1[n*9+(16*C+14)],codeword_buf16[n*10+(16*C+14)],codeword_buf15[n*10+(16*C+14)],codeword_buf14[n*10+(16*C+14)],codeword_buf13[n*10+(16*C+14)],codeword_buf12[n*10+(16*C+14)],codeword_buf11[n*10+(16*C+14)],codeword_buf10[n*10+(16*C+14)],codeword_buf9[n*10+(16*C+14)],codeword_buf8[n*10+(16*C+14)],codeword_buf7[n*10+(16*C+14)],codeword_buf6[n*10+(16*C+14)],codeword_buf5[n*10+(16*C+14)],codeword_buf4[n*10+(16*C+14)],codeword_buf3[n*10+(16*C+14)],codeword_buf2[n*10+(16*C+14)],codeword_buf1[n*10+(16*C+14)],codeword_buf16[n*11+(16*C+14)],codeword_buf15[n*11+(16*C+14)],codeword_buf14[n*11+(16*C+14)],codeword_buf13[n*11+(16*C+14)],codeword_buf12[n*11+(16*C+14)],codeword_buf11[n*11+(16*C+14)],codeword_buf10[n*11+(16*C+14)],codeword_buf9[n*11+(16*C+14)],codeword_buf8[n*11+(16*C+14)],codeword_buf7[n*11+(16*C+14)],codeword_buf6[n*11+(16*C+14)],codeword_buf5[n*11+(16*C+14)],codeword_buf4[n*11+(16*C+14)],codeword_buf3[n*11+(16*C+14)],codeword_buf2[n*11+(16*C+14)],codeword_buf1[n*11+(16*C+14)],codeword_buf16[n*12+(16*C+14)],codeword_buf15[n*12+(16*C+14)],codeword_buf14[n*12+(16*C+14)],codeword_buf13[n*12+(16*C+14)],codeword_buf12[n*12+(16*C+14)],codeword_buf11[n*12+(16*C+14)],codeword_buf10[n*12+(16*C+14)],codeword_buf9[n*12+(16*C+14)],codeword_buf8[n*12+(16*C+14)],codeword_buf7[n*12+(16*C+14)],codeword_buf6[n*12+(16*C+14)],codeword_buf5[n*12+(16*C+14)],codeword_buf4[n*12+(16*C+14)],codeword_buf3[n*12+(16*C+14)],codeword_buf2[n*12+(16*C+14)],codeword_buf1[n*12+(16*C+14)],codeword_buf16[n*13+(16*C+14)],codeword_buf15[n*13+(16*C+14)],codeword_buf14[n*13+(16*C+14)],codeword_buf13[n*13+(16*C+14)],codeword_buf12[n*13+(16*C+14)],codeword_buf11[n*13+(16*C+14)],codeword_buf10[n*13+(16*C+14)],codeword_buf9[n*13+(16*C+14)],codeword_buf8[n*13+(16*C+14)],codeword_buf7[n*13+(16*C+14)],codeword_buf6[n*13+(16*C+14)],codeword_buf5[n*13+(16*C+14)],codeword_buf4[n*13+(16*C+14)],codeword_buf3[n*13+(16*C+14)],codeword_buf2[n*13+(16*C+14)],codeword_buf1[n*13+(16*C+14)],codeword_buf16[n*14+(16*C+14)],codeword_buf15[n*14+(16*C+14)],codeword_buf14[n*14+(16*C+14)],codeword_buf13[n*14+(16*C+14)],codeword_buf12[n*14+(16*C+14)],codeword_buf11[n*14+(16*C+14)],codeword_buf10[n*14+(16*C+14)],codeword_buf9[n*14+(16*C+14)],codeword_buf8[n*14+(16*C+14)],codeword_buf7[n*14+(16*C+14)],codeword_buf6[n*14+(16*C+14)],codeword_buf5[n*14+(16*C+14)],codeword_buf4[n*14+(16*C+14)],codeword_buf3[n*14+(16*C+14)],codeword_buf2[n*14+(16*C+14)],codeword_buf1[n*14+(16*C+14)],codeword_buf16[n*15+(16*C+14)],codeword_buf15[n*15+(16*C+14)],codeword_buf14[n*15+(16*C+14)],codeword_buf13[n*15+(16*C+14)],codeword_buf12[n*15+(16*C+14)],codeword_buf11[n*15+(16*C+14)],codeword_buf10[n*15+(16*C+14)],codeword_buf9[n*15+(16*C+14)],codeword_buf8[n*15+(16*C+14)],codeword_buf7[n*15+(16*C+14)],codeword_buf6[n*15+(16*C+14)],codeword_buf5[n*15+(16*C+14)],codeword_buf4[n*15+(16*C+14)],codeword_buf3[n*15+(16*C+14)],codeword_buf2[n*15+(16*C+14)],codeword_buf1[n*15+(16*C+14)]};
                            in_rec16 <= {codeword_buf16[n*0+(16*C+15)],codeword_buf15[n*0+(16*C+15)],codeword_buf14[n*0+(16*C+15)],codeword_buf13[n*0+(16*C+15)],codeword_buf12[n*0+(16*C+15)],codeword_buf11[n*0+(16*C+15)],codeword_buf10[n*0+(16*C+15)],codeword_buf9[n*0+(16*C+15)],codeword_buf8[n*0+(16*C+15)],codeword_buf7[n*0+(16*C+15)],codeword_buf6[n*0+(16*C+15)],codeword_buf5[n*0+(16*C+15)],codeword_buf4[n*0+(16*C+15)],codeword_buf3[n*0+(16*C+15)],codeword_buf2[n*0+(16*C+15)],codeword_buf1[n*0+(16*C+15)],codeword_buf16[n*1+(16*C+15)],codeword_buf15[n*1+(16*C+15)],codeword_buf14[n*1+(16*C+15)],codeword_buf13[n*1+(16*C+15)],codeword_buf12[n*1+(16*C+15)],codeword_buf11[n*1+(16*C+15)],codeword_buf10[n*1+(16*C+15)],codeword_buf9[n*1+(16*C+15)],codeword_buf8[n*1+(16*C+15)],codeword_buf7[n*1+(16*C+15)],codeword_buf6[n*1+(16*C+15)],codeword_buf5[n*1+(16*C+15)],codeword_buf4[n*1+(16*C+15)],codeword_buf3[n*1+(16*C+15)],codeword_buf2[n*1+(16*C+15)],codeword_buf1[n*1+(16*C+15)],codeword_buf16[n*2+(16*C+15)],codeword_buf15[n*2+(16*C+15)],codeword_buf14[n*2+(16*C+15)],codeword_buf13[n*2+(16*C+15)],codeword_buf12[n*2+(16*C+15)],codeword_buf11[n*2+(16*C+15)],codeword_buf10[n*2+(16*C+15)],codeword_buf9[n*2+(16*C+15)],codeword_buf8[n*2+(16*C+15)],codeword_buf7[n*2+(16*C+15)],codeword_buf6[n*2+(16*C+15)],codeword_buf5[n*2+(16*C+15)],codeword_buf4[n*2+(16*C+15)],codeword_buf3[n*2+(16*C+15)],codeword_buf2[n*2+(16*C+15)],codeword_buf1[n*2+(16*C+15)],codeword_buf16[n*3+(16*C+15)],codeword_buf15[n*3+(16*C+15)],codeword_buf14[n*3+(16*C+15)],codeword_buf13[n*3+(16*C+15)],codeword_buf12[n*3+(16*C+15)],codeword_buf11[n*3+(16*C+15)],codeword_buf10[n*3+(16*C+15)],codeword_buf9[n*3+(16*C+15)],codeword_buf8[n*3+(16*C+15)],codeword_buf7[n*3+(16*C+15)],codeword_buf6[n*3+(16*C+15)],codeword_buf5[n*3+(16*C+15)],codeword_buf4[n*3+(16*C+15)],codeword_buf3[n*3+(16*C+15)],codeword_buf2[n*3+(16*C+15)],codeword_buf1[n*3+(16*C+15)],codeword_buf16[n*4+(16*C+15)],codeword_buf15[n*4+(16*C+15)],codeword_buf14[n*4+(16*C+15)],codeword_buf13[n*4+(16*C+15)],codeword_buf12[n*4+(16*C+15)],codeword_buf11[n*4+(16*C+15)],codeword_buf10[n*4+(16*C+15)],codeword_buf9[n*4+(16*C+15)],codeword_buf8[n*4+(16*C+15)],codeword_buf7[n*4+(16*C+15)],codeword_buf6[n*4+(16*C+15)],codeword_buf5[n*4+(16*C+15)],codeword_buf4[n*4+(16*C+15)],codeword_buf3[n*4+(16*C+15)],codeword_buf2[n*4+(16*C+15)],codeword_buf1[n*4+(16*C+15)],codeword_buf16[n*5+(16*C+15)],codeword_buf15[n*5+(16*C+15)],codeword_buf14[n*5+(16*C+15)],codeword_buf13[n*5+(16*C+15)],codeword_buf12[n*5+(16*C+15)],codeword_buf11[n*5+(16*C+15)],codeword_buf10[n*5+(16*C+15)],codeword_buf9[n*5+(16*C+15)],codeword_buf8[n*5+(16*C+15)],codeword_buf7[n*5+(16*C+15)],codeword_buf6[n*5+(16*C+15)],codeword_buf5[n*5+(16*C+15)],codeword_buf4[n*5+(16*C+15)],codeword_buf3[n*5+(16*C+15)],codeword_buf2[n*5+(16*C+15)],codeword_buf1[n*5+(16*C+15)],codeword_buf16[n*6+(16*C+15)],codeword_buf15[n*6+(16*C+15)],codeword_buf14[n*6+(16*C+15)],codeword_buf13[n*6+(16*C+15)],codeword_buf12[n*6+(16*C+15)],codeword_buf11[n*6+(16*C+15)],codeword_buf10[n*6+(16*C+15)],codeword_buf9[n*6+(16*C+15)],codeword_buf8[n*6+(16*C+15)],codeword_buf7[n*6+(16*C+15)],codeword_buf6[n*6+(16*C+15)],codeword_buf5[n*6+(16*C+15)],codeword_buf4[n*6+(16*C+15)],codeword_buf3[n*6+(16*C+15)],codeword_buf2[n*6+(16*C+15)],codeword_buf1[n*6+(16*C+15)],codeword_buf16[n*7+(16*C+15)],codeword_buf15[n*7+(16*C+15)],codeword_buf14[n*7+(16*C+15)],codeword_buf13[n*7+(16*C+15)],codeword_buf12[n*7+(16*C+15)],codeword_buf11[n*7+(16*C+15)],codeword_buf10[n*7+(16*C+15)],codeword_buf9[n*7+(16*C+15)],codeword_buf8[n*7+(16*C+15)],codeword_buf7[n*7+(16*C+15)],codeword_buf6[n*7+(16*C+15)],codeword_buf5[n*7+(16*C+15)],codeword_buf4[n*7+(16*C+15)],codeword_buf3[n*7+(16*C+15)],codeword_buf2[n*7+(16*C+15)],codeword_buf1[n*7+(16*C+15)],codeword_buf16[n*8+(16*C+15)],codeword_buf15[n*8+(16*C+15)],codeword_buf14[n*8+(16*C+15)],codeword_buf13[n*8+(16*C+15)],codeword_buf12[n*8+(16*C+15)],codeword_buf11[n*8+(16*C+15)],codeword_buf10[n*8+(16*C+15)],codeword_buf9[n*8+(16*C+15)],codeword_buf8[n*8+(16*C+15)],codeword_buf7[n*8+(16*C+15)],codeword_buf6[n*8+(16*C+15)],codeword_buf5[n*8+(16*C+15)],codeword_buf4[n*8+(16*C+15)],codeword_buf3[n*8+(16*C+15)],codeword_buf2[n*8+(16*C+15)],codeword_buf1[n*8+(16*C+15)],codeword_buf16[n*9+(16*C+15)],codeword_buf15[n*9+(16*C+15)],codeword_buf14[n*9+(16*C+15)],codeword_buf13[n*9+(16*C+15)],codeword_buf12[n*9+(16*C+15)],codeword_buf11[n*9+(16*C+15)],codeword_buf10[n*9+(16*C+15)],codeword_buf9[n*9+(16*C+15)],codeword_buf8[n*9+(16*C+15)],codeword_buf7[n*9+(16*C+15)],codeword_buf6[n*9+(16*C+15)],codeword_buf5[n*9+(16*C+15)],codeword_buf4[n*9+(16*C+15)],codeword_buf3[n*9+(16*C+15)],codeword_buf2[n*9+(16*C+15)],codeword_buf1[n*9+(16*C+15)],codeword_buf16[n*10+(16*C+15)],codeword_buf15[n*10+(16*C+15)],codeword_buf14[n*10+(16*C+15)],codeword_buf13[n*10+(16*C+15)],codeword_buf12[n*10+(16*C+15)],codeword_buf11[n*10+(16*C+15)],codeword_buf10[n*10+(16*C+15)],codeword_buf9[n*10+(16*C+15)],codeword_buf8[n*10+(16*C+15)],codeword_buf7[n*10+(16*C+15)],codeword_buf6[n*10+(16*C+15)],codeword_buf5[n*10+(16*C+15)],codeword_buf4[n*10+(16*C+15)],codeword_buf3[n*10+(16*C+15)],codeword_buf2[n*10+(16*C+15)],codeword_buf1[n*10+(16*C+15)],codeword_buf16[n*11+(16*C+15)],codeword_buf15[n*11+(16*C+15)],codeword_buf14[n*11+(16*C+15)],codeword_buf13[n*11+(16*C+15)],codeword_buf12[n*11+(16*C+15)],codeword_buf11[n*11+(16*C+15)],codeword_buf10[n*11+(16*C+15)],codeword_buf9[n*11+(16*C+15)],codeword_buf8[n*11+(16*C+15)],codeword_buf7[n*11+(16*C+15)],codeword_buf6[n*11+(16*C+15)],codeword_buf5[n*11+(16*C+15)],codeword_buf4[n*11+(16*C+15)],codeword_buf3[n*11+(16*C+15)],codeword_buf2[n*11+(16*C+15)],codeword_buf1[n*11+(16*C+15)],codeword_buf16[n*12+(16*C+15)],codeword_buf15[n*12+(16*C+15)],codeword_buf14[n*12+(16*C+15)],codeword_buf13[n*12+(16*C+15)],codeword_buf12[n*12+(16*C+15)],codeword_buf11[n*12+(16*C+15)],codeword_buf10[n*12+(16*C+15)],codeword_buf9[n*12+(16*C+15)],codeword_buf8[n*12+(16*C+15)],codeword_buf7[n*12+(16*C+15)],codeword_buf6[n*12+(16*C+15)],codeword_buf5[n*12+(16*C+15)],codeword_buf4[n*12+(16*C+15)],codeword_buf3[n*12+(16*C+15)],codeword_buf2[n*12+(16*C+15)],codeword_buf1[n*12+(16*C+15)],codeword_buf16[n*13+(16*C+15)],codeword_buf15[n*13+(16*C+15)],codeword_buf14[n*13+(16*C+15)],codeword_buf13[n*13+(16*C+15)],codeword_buf12[n*13+(16*C+15)],codeword_buf11[n*13+(16*C+15)],codeword_buf10[n*13+(16*C+15)],codeword_buf9[n*13+(16*C+15)],codeword_buf8[n*13+(16*C+15)],codeword_buf7[n*13+(16*C+15)],codeword_buf6[n*13+(16*C+15)],codeword_buf5[n*13+(16*C+15)],codeword_buf4[n*13+(16*C+15)],codeword_buf3[n*13+(16*C+15)],codeword_buf2[n*13+(16*C+15)],codeword_buf1[n*13+(16*C+15)],codeword_buf16[n*14+(16*C+15)],codeword_buf15[n*14+(16*C+15)],codeword_buf14[n*14+(16*C+15)],codeword_buf13[n*14+(16*C+15)],codeword_buf12[n*14+(16*C+15)],codeword_buf11[n*14+(16*C+15)],codeword_buf10[n*14+(16*C+15)],codeword_buf9[n*14+(16*C+15)],codeword_buf8[n*14+(16*C+15)],codeword_buf7[n*14+(16*C+15)],codeword_buf6[n*14+(16*C+15)],codeword_buf5[n*14+(16*C+15)],codeword_buf4[n*14+(16*C+15)],codeword_buf3[n*14+(16*C+15)],codeword_buf2[n*14+(16*C+15)],codeword_buf1[n*14+(16*C+15)],codeword_buf16[n*15+(16*C+15)],codeword_buf15[n*15+(16*C+15)],codeword_buf14[n*15+(16*C+15)],codeword_buf13[n*15+(16*C+15)],codeword_buf12[n*15+(16*C+15)],codeword_buf11[n*15+(16*C+15)],codeword_buf10[n*15+(16*C+15)],codeword_buf9[n*15+(16*C+15)],codeword_buf8[n*15+(16*C+15)],codeword_buf7[n*15+(16*C+15)],codeword_buf6[n*15+(16*C+15)],codeword_buf5[n*15+(16*C+15)],codeword_buf4[n*15+(16*C+15)],codeword_buf3[n*15+(16*C+15)],codeword_buf2[n*15+(16*C+15)],codeword_buf1[n*15+(16*C+15)]};
    
                        
                            C <= C + 1;     // Decrease the C value
                        end
                        
                        // Shift the buffer values to save the new column decoded values
                        codeword_buf2_1  <= (codeword_buf2_1  << n);
                        codeword_buf2_2  <= (codeword_buf2_2  << n);
                        codeword_buf2_3  <= (codeword_buf2_3  << n);
                        codeword_buf2_4  <= (codeword_buf2_4  << n);
                        codeword_buf2_5  <= (codeword_buf2_5  << n);
                        codeword_buf2_6  <= (codeword_buf2_6  << n);
                        codeword_buf2_7  <= (codeword_buf2_7  << n);
                        codeword_buf2_8  <= (codeword_buf2_8  << n);
                        codeword_buf2_9  <= (codeword_buf2_9  << n);
                        codeword_buf2_10 <= (codeword_buf2_10 << n);
                        codeword_buf2_11 <= (codeword_buf2_11 << n);
                        codeword_buf2_12 <= (codeword_buf2_12 << n);
                        codeword_buf2_13 <= (codeword_buf2_13 << n);
                        codeword_buf2_14 <= (codeword_buf2_14 << n);
                        codeword_buf2_15 <= (codeword_buf2_15 << n);
                        codeword_buf2_16 <= (codeword_buf2_16 << n);
                        
                        // Save the column decoded values in the buffer
                        codeword_buf2_1[(n-1):0]  <= out_dec1;
                        codeword_buf2_2[(n-1):0]  <= out_dec2;
                        codeword_buf2_3[(n-1):0]  <= out_dec3;
                        codeword_buf2_4[(n-1):0]  <= out_dec4;
                        codeword_buf2_5[(n-1):0]  <= out_dec5;
                        codeword_buf2_6[(n-1):0]  <= out_dec6;
                        codeword_buf2_7[(n-1):0]  <= out_dec7;
                        codeword_buf2_8[(n-1):0]  <= out_dec8;
                        codeword_buf2_9[(n-1):0]  <= out_dec9;
                        codeword_buf2_10[(n-1):0] <= out_dec10;
                        codeword_buf2_11[(n-1):0] <= out_dec11;
                        codeword_buf2_12[(n-1):0] <= out_dec12;
                        codeword_buf2_13[(n-1):0] <= out_dec13;
                        codeword_buf2_14[(n-1):0] <= out_dec14;
                        codeword_buf2_15[(n-1):0] <= out_dec15;
                        codeword_buf2_16[(n-1):0] <= out_dec16;
                        
    //                    if (counter == 4'h8)
    //                        valid1 <= 1'b1;
    //                    else
    
                        valid1 <= 1'b0;
                        
                        // Change the valid2 values to inform the datapath, that the decoded codewords are valid
                        if ((counter >= 6'd30)&&(counter < 6'd45))
                            valid2 <= 1'b1;
                        else
                            valid2 <= 1'b0;
                            
//                        if (counter == 6'd45)
//                            valid_err <= 1'b0;
//                        else 
//                            valid_err <= 1'b0;
                        
                        // If the counter is in this range output the assigned values to the registers, else assign x
                        if ((counter > 6'd29)&&(rounds == 1)) begin
                            dec1  <= out_dec1;
                            dec2  <= out_dec2;
                            dec3  <= out_dec3;
                            dec4  <= out_dec4;
                            dec5  <= out_dec5;
                            dec6  <= out_dec6;
                            dec7  <= out_dec7;
                            dec8  <= out_dec8;
                            dec9  <= out_dec9;
                            dec10 <= out_dec10;
                            dec11 <= out_dec11;
                            dec12 <= out_dec12;
                            dec13 <= out_dec13;
                            dec14 <= out_dec14;
                            dec15 <= out_dec15;
                            dec16 <= out_dec16;
                        end else begin
                            dec1  <= 256'bx;
                            dec2  <= 256'bx;
                            dec3  <= 256'bx;
                            dec4  <= 256'bx;
                            dec5  <= 256'bx;
                            dec6  <= 256'bx;
                            dec7  <= 256'bx;
                            dec8  <= 256'bx;
                            dec9  <= 256'bx;
                            dec10 <= 256'bx;
                            dec11 <= 256'bx;
                            dec12 <= 256'bx;
                            dec13 <= 256'bx;
                            dec14 <= 256'bx;
                            dec15 <= 256'bx;
                            dec16 <= 256'bx;
                        end
                        
    //                    // If the counter value is more than or equal to 41, send the signal to start encoding
    //                    if (counter >= 6'd42)
    //                        hold_enc <= 1'b1;
    //                    else
    //                        hold_enc <= 1'b0;
                        
                        // Change the counter value and rounds value accordingly
                        if (counter < 6'd50)
                            counter <= counter + 4'b1;
                        else if ((counter == 6'd50)&&(rounds > 1)) begin
                            counter <= 6'd23; 
                            rounds <= rounds - 1;
                        end else begin
                            counter <= 4'b0;
                            rounds <= iter * 2;
                            C <= 4'd0;
                        end
                        
                    end else begin
                    
                        if (counter == 6'd46)
                            valid_err <= 1'b1;
                        else 
                            valid_err <= 1'b0;
                    
                        if (counter < 6'd50)
                            counter <= counter + 4'b1;
                        else if ((counter == 6'd50)&&(rounds > 1)) begin
                            counter <= 6'd23; 
                            rounds <= rounds - 1;
                        end else begin
                            counter <= 4'b0;
                            rounds <= iter * 2;
                            C <= 4'd0;
                        end
                        
                        valid2 <= 1'b0;
                    end
                end
                //// End of the column decoding block ////
            end
            //// End of the decoding ////
        
        // If the system is OFF       
        end else begin
            counter <= 4'b0;
            hold <= 1'b0;
            valid1 <= 1'b0;
            valid2 <= 1'b0;
            rounds <= iter*2;
            hold_enc <= 1'b1;
            C <= 4'd0;
        end
    end
        
endmodule
