`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/13/2024 02:57:45 PM
// Design Name: 
// Module Name: interleaver_128
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module interleaver_2048(
    input clk,
    input reset,
    input wire [4095:0] in,
    output reg [4095:0] out
    );

    always @(posedge clk) begin
        out[0] <= in[1937]; 
        out[1] <= in[2448]; 
        out[2] <= in[1755]; 
        out[3] <= in[3464]; 
        out[4] <= in[993]; 
        out[5] <= in[2232]; 
        out[6] <= in[1244]; 
        out[7] <= in[3]; 
        out[8] <= in[3974]; 
        out[9] <= in[1676]; 
        out[10] <= in[4016]; 
        out[11] <= in[1356]; 
        out[12] <= in[753]; 
        out[13] <= in[3624]; 
        out[14] <= in[487]; 
        out[15] <= in[3268]; 
        out[16] <= in[370]; 
        out[17] <= in[1349]; 
        out[18] <= in[2578]; 
        out[19] <= in[1129]; 
        out[20] <= in[1173]; 
        out[21] <= in[2925]; 
        out[22] <= in[1493]; 
        out[23] <= in[3727]; 
        out[24] <= in[2314]; 
        out[25] <= in[2575]; 
        out[26] <= in[1990]; 
        out[27] <= in[2096]; 
        out[28] <= in[2704]; 
        out[29] <= in[520]; 
        out[30] <= in[1801]; 
        out[31] <= in[1727]; 
        out[32] <= in[2752]; 
        out[33] <= in[1759]; 
        out[34] <= in[2963]; 
        out[35] <= in[2868]; 
        out[36] <= in[2642]; 
        out[37] <= in[2551]; 
        out[38] <= in[525]; 
        out[39] <= in[203]; 
        out[40] <= in[682]; 
        out[41] <= in[1882]; 
        out[42] <= in[3500]; 
        out[43] <= in[4028]; 
        out[44] <= in[3220]; 
        out[45] <= in[113]; 
        out[46] <= in[2479]; 
        out[47] <= in[999]; 
        out[48] <= in[1768]; 
        out[49] <= in[2184]; 
        out[50] <= in[3489]; 
        out[51] <= in[2533]; 
        out[52] <= in[3385]; 
        out[53] <= in[1262]; 
        out[54] <= in[355]; 
        out[55] <= in[2385]; 
        out[56] <= in[3139]; 
        out[57] <= in[931]; 
        out[58] <= in[2259]; 
        out[59] <= in[2745]; 
        out[60] <= in[2847]; 
        out[61] <= in[3713]; 
        out[62] <= in[1729]; 
        out[63] <= in[1604]; 
        out[64] <= in[563]; 
        out[65] <= in[3336]; 
        out[66] <= in[2010]; 
        out[67] <= in[3947]; 
        out[68] <= in[236]; 
        out[69] <= in[30]; 
        out[70] <= in[2214]; 
        out[71] <= in[2703]; 
        out[72] <= in[3081]; 
        out[73] <= in[1248]; 
        out[74] <= in[484]; 
        out[75] <= in[3509]; 
        out[76] <= in[107]; 
        out[77] <= in[2702]; 
        out[78] <= in[2565]; 
        out[79] <= in[3032]; 
        out[80] <= in[1706]; 
        out[81] <= in[1847]; 
        out[82] <= in[2222]; 
        out[83] <= in[2759]; 
        out[84] <= in[512]; 
        out[85] <= in[2472]; 
        out[86] <= in[1997]; 
        out[87] <= in[1589]; 
        out[88] <= in[3894]; 
        out[89] <= in[1996]; 
        out[90] <= in[199]; 
        out[91] <= in[3843]; 
        out[92] <= in[2646]; 
        out[93] <= in[1459]; 
        out[94] <= in[1892]; 
        out[95] <= in[2645]; 
        out[96] <= in[4051]; 
        out[97] <= in[1597]; 
        out[98] <= in[2741]; 
        out[99] <= in[1235]; 
        out[100] <= in[647]; 
        out[101] <= in[2373]; 
        out[102] <= in[1329]; 
        out[103] <= in[260]; 
        out[104] <= in[3225]; 
        out[105] <= in[275]; 
        out[106] <= in[3942]; 
        out[107] <= in[3473]; 
        out[108] <= in[1764]; 
        out[109] <= in[2522]; 
        out[110] <= in[293]; 
        out[111] <= in[3794]; 
        out[112] <= in[1295]; 
        out[113] <= in[1399]; 
        out[114] <= in[412]; 
        out[115] <= in[969]; 
        out[116] <= in[2927]; 
        out[117] <= in[2885]; 
        out[118] <= in[1778]; 
        out[119] <= in[2310]; 
        out[120] <= in[2527]; 
        out[121] <= in[1974]; 
        out[122] <= in[2248]; 
        out[123] <= in[2996]; 
        out[124] <= in[2306]; 
        out[125] <= in[3479]; 
        out[126] <= in[31]; 
        out[127] <= in[3371]; 
        out[128] <= in[2371]; 
        out[129] <= in[3536]; 
        out[130] <= in[2604]; 
        out[131] <= in[252]; 
        out[132] <= in[3575]; 
        out[133] <= in[3253]; 
        out[134] <= in[205]; 
        out[135] <= in[1450]; 
        out[136] <= in[3282]; 
        out[137] <= in[3392]; 
        out[138] <= in[1328]; 
        out[139] <= in[2104]; 
        out[140] <= in[1134]; 
        out[141] <= in[530]; 
        out[142] <= in[2517]; 
        out[143] <= in[1814]; 
        out[144] <= in[1398]; 
        out[145] <= in[3349]; 
        out[146] <= in[2554]; 
        out[147] <= in[3660]; 
        out[148] <= in[3332]; 
        out[149] <= in[155]; 
        out[150] <= in[102]; 
        out[151] <= in[619]; 
        out[152] <= in[1157]; 
        out[153] <= in[2713]; 
        out[154] <= in[3643]; 
        out[155] <= in[2224]; 
        out[156] <= in[378]; 
        out[157] <= in[3816]; 
        out[158] <= in[1461]; 
        out[159] <= in[948]; 
        out[160] <= in[1647]; 
        out[161] <= in[3102]; 
        out[162] <= in[2419]; 
        out[163] <= in[167]; 
        out[164] <= in[1723]; 
        out[165] <= in[367]; 
        out[166] <= in[1347]; 
        out[167] <= in[1746]; 
        out[168] <= in[609]; 
        out[169] <= in[1439]; 
        out[170] <= in[3465]; 
        out[171] <= in[2296]; 
        out[172] <= in[2663]; 
        out[173] <= in[861]; 
        out[174] <= in[2539]; 
        out[175] <= in[2454]; 
        out[176] <= in[122]; 
        out[177] <= in[3683]; 
        out[178] <= in[3034]; 
        out[179] <= in[2907]; 
        out[180] <= in[980]; 
        out[181] <= in[1799]; 
        out[182] <= in[2157]; 
        out[183] <= in[1374]; 
        out[184] <= in[1179]; 
        out[185] <= in[1204]; 
        out[186] <= in[2499]; 
        out[187] <= in[627]; 
        out[188] <= in[2732]; 
        out[189] <= in[3384]; 
        out[190] <= in[1958]; 
        out[191] <= in[52]; 
        out[192] <= in[50]; 
        out[193] <= in[499]; 
        out[194] <= in[543]; 
        out[195] <= in[2758]; 
        out[196] <= in[1857]; 
        out[197] <= in[1805]; 
        out[198] <= in[2431]; 
        out[199] <= in[2696]; 
        out[200] <= in[4044]; 
        out[201] <= in[2507]; 
        out[202] <= in[2046]; 
        out[203] <= in[3918]; 
        out[204] <= in[3127]; 
        out[205] <= in[1740]; 
        out[206] <= in[3451]; 
        out[207] <= in[3983]; 
        out[208] <= in[1054]; 
        out[209] <= in[1327]; 
        out[210] <= in[2666]; 
        out[211] <= in[2570]; 
        out[212] <= in[2156]; 
        out[213] <= in[3052]; 
        out[214] <= in[3140]; 
        out[215] <= in[1691]; 
        out[216] <= in[290]; 
        out[217] <= in[705]; 
        out[218] <= in[574]; 
        out[219] <= in[1476]; 
        out[220] <= in[3966]; 
        out[221] <= in[828]; 
        out[222] <= in[1786]; 
        out[223] <= in[2223]; 
        out[224] <= in[2105]; 
        out[225] <= in[3166]; 
        out[226] <= in[1619]; 
        out[227] <= in[1842]; 
        out[228] <= in[1827]; 
        out[229] <= in[1107]; 
        out[230] <= in[3825]; 
        out[231] <= in[2583]; 
        out[232] <= in[1481]; 
        out[233] <= in[3414]; 
        out[234] <= in[2960]; 
        out[235] <= in[532]; 
        out[236] <= in[3099]; 
        out[237] <= in[1562]; 
        out[238] <= in[3357]; 
        out[239] <= in[3805]; 
        out[240] <= in[838]; 
        out[241] <= in[1655]; 
        out[242] <= in[1737]; 
        out[243] <= in[1927]; 
        out[244] <= in[982]; 
        out[245] <= in[3141]; 
        out[246] <= in[1670]; 
        out[247] <= in[4023]; 
        out[248] <= in[3310]; 
        out[249] <= in[3897]; 
        out[250] <= in[2075]; 
        out[251] <= in[871]; 
        out[252] <= in[3405]; 
        out[253] <= in[2012]; 
        out[254] <= in[2086]; 
        out[255] <= in[765]; 
        out[256] <= in[380]; 
        out[257] <= in[939]; 
        out[258] <= in[3776]; 
        out[259] <= in[3513]; 
        out[260] <= in[1550]; 
        out[261] <= in[1361]; 
        out[262] <= in[3952]; 
        out[263] <= in[2633]; 
        out[264] <= in[3173]; 
        out[265] <= in[1028]; 
        out[266] <= in[1339]; 
        out[267] <= in[2611]; 
        out[268] <= in[2335]; 
        out[269] <= in[1806]; 
        out[270] <= in[2069]; 
        out[271] <= in[3296]; 
        out[272] <= in[938]; 
        out[273] <= in[3186]; 
        out[274] <= in[446]; 
        out[275] <= in[851]; 
        out[276] <= in[2797]; 
        out[277] <= in[3468]; 
        out[278] <= in[746]; 
        out[279] <= in[3766]; 
        out[280] <= in[3540]; 
        out[281] <= in[2355]; 
        out[282] <= in[1823]; 
        out[283] <= in[3056]; 
        out[284] <= in[3302]; 
        out[285] <= in[1658]; 
        out[286] <= in[3292]; 
        out[287] <= in[2846]; 
        out[288] <= in[395]; 
        out[289] <= in[1279]; 
        out[290] <= in[1519]; 
        out[291] <= in[604]; 
        out[292] <= in[1158]; 
        out[293] <= in[2682]; 
        out[294] <= in[2816]; 
        out[295] <= in[2257]; 
        out[296] <= in[569]; 
        out[297] <= in[1689]; 
        out[298] <= in[3343]; 
        out[299] <= in[896]; 
        out[300] <= in[1736]; 
        out[301] <= in[2070]; 
        out[302] <= in[2970]; 
        out[303] <= in[3162]; 
        out[304] <= in[1128]; 
        out[305] <= in[3557]; 
        out[306] <= in[3745]; 
        out[307] <= in[119]; 
        out[308] <= in[3433]; 
        out[309] <= in[2841]; 
        out[310] <= in[4081]; 
        out[311] <= in[3986]; 
        out[312] <= in[1355]; 
        out[313] <= in[3854]; 
        out[314] <= in[3375]; 
        out[315] <= in[3158]; 
        out[316] <= in[1633]; 
        out[317] <= in[2928]; 
        out[318] <= in[2665]; 
        out[319] <= in[1527]; 
        out[320] <= in[4010]; 
        out[321] <= in[2924]; 
        out[322] <= in[4076]; 
        out[323] <= in[2017]; 
        out[324] <= in[400]; 
        out[325] <= in[3633]; 
        out[326] <= in[3168]; 
        out[327] <= in[3101]; 
        out[328] <= in[1207]; 
        out[329] <= in[129]; 
        out[330] <= in[1953]; 
        out[331] <= in[1052]; 
        out[332] <= in[975]; 
        out[333] <= in[4009]; 
        out[334] <= in[1039]; 
        out[335] <= in[928]; 
        out[336] <= in[3378]; 
        out[337] <= in[2946]; 
        out[338] <= in[3243]; 
        out[339] <= in[1626]; 
        out[340] <= in[2993]; 
        out[341] <= in[1893]; 
        out[342] <= in[1475]; 
        out[343] <= in[2258]; 
        out[344] <= in[2410]; 
        out[345] <= in[51]; 
        out[346] <= in[1288]; 
        out[347] <= in[1686]; 
        out[348] <= in[2150]; 
        out[349] <= in[2931]; 
        out[350] <= in[2973]; 
        out[351] <= in[2897]; 
        out[352] <= in[2364]; 
        out[353] <= in[2941]; 
        out[354] <= in[1187]; 
        out[355] <= in[1930]; 
        out[356] <= in[2675]; 
        out[357] <= in[3115]; 
        out[358] <= in[278]; 
        out[359] <= in[2894]; 
        out[360] <= in[2524]; 
        out[361] <= in[981]; 
        out[362] <= in[3364]; 
        out[363] <= in[3437]; 
        out[364] <= in[3690]; 
        out[365] <= in[924]; 
        out[366] <= in[3287]; 
        out[367] <= in[509]; 
        out[368] <= in[3033]; 
        out[369] <= in[185]; 
        out[370] <= in[1600]; 
        out[371] <= in[2923]; 
        out[372] <= in[2451]; 
        out[373] <= in[1609]; 
        out[374] <= in[3455]; 
        out[375] <= in[777]; 
        out[376] <= in[2720]; 
        out[377] <= in[811]; 
        out[378] <= in[1404]; 
        out[379] <= in[1079]; 
        out[380] <= in[1971]; 
        out[381] <= in[2395]; 
        out[382] <= in[3886]; 
        out[383] <= in[3320]; 
        out[384] <= in[2095]; 
        out[385] <= in[3757]; 
        out[386] <= in[1023]; 
        out[387] <= in[3929]; 
        out[388] <= in[3953]; 
        out[389] <= in[2831]; 
        out[390] <= in[3807]; 
        out[391] <= in[3178]; 
        out[392] <= in[1744]; 
        out[393] <= in[25]; 
        out[394] <= in[4032]; 
        out[395] <= in[1767]; 
        out[396] <= in[1675]; 
        out[397] <= in[2975]; 
        out[398] <= in[1710]; 
        out[399] <= in[3553]; 
        out[400] <= in[2485]; 
        out[401] <= in[3635]; 
        out[402] <= in[951]; 
        out[403] <= in[3070]; 
        out[404] <= in[4043]; 
        out[405] <= in[1153]; 
        out[406] <= in[799]; 
        out[407] <= in[3872]; 
        out[408] <= in[2980]; 
        out[409] <= in[1379]; 
        out[410] <= in[388]; 
        out[411] <= in[3839]; 
        out[412] <= in[1742]; 
        out[413] <= in[1918]; 
        out[414] <= in[1409]; 
        out[415] <= in[1165]; 
        out[416] <= in[2346]; 
        out[417] <= in[1067]; 
        out[418] <= in[3985]; 
        out[419] <= in[3169]; 
        out[420] <= in[3211]; 
        out[421] <= in[3359]; 
        out[422] <= in[990]; 
        out[423] <= in[1097]; 
        out[424] <= in[246]; 
        out[425] <= in[3855]; 
        out[426] <= in[966]; 
        out[427] <= in[3480]; 
        out[428] <= in[463]; 
        out[429] <= in[152]; 
        out[430] <= in[2986]; 
        out[431] <= in[3949]; 
        out[432] <= in[1784]; 
        out[433] <= in[3779]; 
        out[434] <= in[2241]; 
        out[435] <= in[3959]; 
        out[436] <= in[2538]; 
        out[437] <= in[3712]; 
        out[438] <= in[1045]; 
        out[439] <= in[2060]; 
        out[440] <= in[2350]; 
        out[441] <= in[174]; 
        out[442] <= in[1919]; 
        out[443] <= in[114]; 
        out[444] <= in[1564]; 
        out[445] <= in[3400]; 
        out[446] <= in[2458]; 
        out[447] <= in[1557]; 
        out[448] <= in[3891]; 
        out[449] <= in[1256]; 
        out[450] <= in[1215]; 
        out[451] <= in[154]; 
        out[452] <= in[492]; 
        out[453] <= in[1512]; 
        out[454] <= in[3814]; 
        out[455] <= in[1280]; 
        out[456] <= in[161]; 
        out[457] <= in[1555]; 
        out[458] <= in[527]; 
        out[459] <= in[1007]; 
        out[460] <= in[769]; 
        out[461] <= in[27]; 
        out[462] <= in[3791]; 
        out[463] <= in[1650]; 
        out[464] <= in[637]; 
        out[465] <= in[3708]; 
        out[466] <= in[3812]; 
        out[467] <= in[2342]; 
        out[468] <= in[2624]; 
        out[469] <= in[654]; 
        out[470] <= in[1278]; 
        out[471] <= in[3116]; 
        out[472] <= in[2730]; 
        out[473] <= in[671]; 
        out[474] <= in[3874]; 
        out[475] <= in[3107]; 
        out[476] <= in[215]; 
        out[477] <= in[3216]; 
        out[478] <= in[1112]; 
        out[479] <= in[2526]; 
        out[480] <= in[3181]; 
        out[481] <= in[3227]; 
        out[482] <= in[3556]; 
        out[483] <= in[1526]; 
        out[484] <= in[140]; 
        out[485] <= in[1998]; 
        out[486] <= in[1147]; 
        out[487] <= in[3134]; 
        out[488] <= in[663]; 
        out[489] <= in[3004]; 
        out[490] <= in[2606]; 
        out[491] <= in[1503]; 
        out[492] <= in[1121]; 
        out[493] <= in[864]; 
        out[494] <= in[3785]; 
        out[495] <= in[3981]; 
        out[496] <= in[703]; 
        out[497] <= in[3058]; 
        out[498] <= in[342]; 
        out[499] <= in[3786]; 
        out[500] <= in[1076]; 
        out[501] <= in[2950]; 
        out[502] <= in[1563]; 
        out[503] <= in[2148]; 
        out[504] <= in[1758]; 
        out[505] <= in[3585]; 
        out[506] <= in[1357]; 
        out[507] <= in[2300]; 
        out[508] <= in[2078]; 
        out[509] <= in[61]; 
        out[510] <= in[1708]; 
        out[511] <= in[796]; 
        out[512] <= in[2810]; 
        out[513] <= in[2299]; 
        out[514] <= in[1160]; 
        out[515] <= in[3103]; 
        out[516] <= in[2515]; 
        out[517] <= in[270]; 
        out[518] <= in[3977]; 
        out[519] <= in[2684]; 
        out[520] <= in[1320]; 
        out[521] <= in[2582]; 
        out[522] <= in[1833]; 
        out[523] <= in[239]; 
        out[524] <= in[1223]; 
        out[525] <= in[729]; 
        out[526] <= in[1632]; 
        out[527] <= in[1267]; 
        out[528] <= in[3482]; 
        out[529] <= in[3999]; 
        out[530] <= in[2026]; 
        out[531] <= in[3212]; 
        out[532] <= in[2028]; 
        out[533] <= in[2509]; 
        out[534] <= in[915]; 
        out[535] <= in[3155]; 
        out[536] <= in[2634]; 
        out[537] <= in[2165]; 
        out[538] <= in[1941]; 
        out[539] <= in[482]; 
        out[540] <= in[441]; 
        out[541] <= in[2734]; 
        out[542] <= in[2376]; 
        out[543] <= in[3495]; 
        out[544] <= in[1995]; 
        out[545] <= in[977]; 
        out[546] <= in[1177]; 
        out[547] <= in[2839]; 
        out[548] <= in[2972]; 
        out[549] <= in[54]; 
        out[550] <= in[3128]; 
        out[551] <= in[3054]; 
        out[552] <= in[1344]; 
        out[553] <= in[2348]; 
        out[554] <= in[2038]; 
        out[555] <= in[2593]; 
        out[556] <= in[1657]; 
        out[557] <= in[3547]; 
        out[558] <= in[2464]; 
        out[559] <= in[2298]; 
        out[560] <= in[3702]; 
        out[561] <= in[3309]; 
        out[562] <= in[1803]; 
        out[563] <= in[1024]; 
        out[564] <= in[164]; 
        out[565] <= in[2892]; 
        out[566] <= in[2261]; 
        out[567] <= in[3501]; 
        out[568] <= in[1794]; 
        out[569] <= in[1698]; 
        out[570] <= in[2307]; 
        out[571] <= in[2881]; 
        out[572] <= in[160]; 
        out[573] <= in[1617]; 
        out[574] <= in[1739]; 
        out[575] <= in[3124]; 
        out[576] <= in[1678]; 
        out[577] <= in[3367]; 
        out[578] <= in[2546]; 
        out[579] <= in[3772]; 
        out[580] <= in[1402]; 
        out[581] <= in[1543]; 
        out[582] <= in[1495]; 
        out[583] <= in[885]; 
        out[584] <= in[1377]; 
        out[585] <= in[1098]; 
        out[586] <= in[3493]; 
        out[587] <= in[419]; 
        out[588] <= in[725]; 
        out[589] <= in[92]; 
        out[590] <= in[3024]; 
        out[591] <= in[1668]; 
        out[592] <= in[4080]; 
        out[593] <= in[1087]; 
        out[594] <= in[3429]; 
        out[595] <= in[551]; 
        out[596] <= in[1588]; 
        out[597] <= in[1321]; 
        out[598] <= in[3300]; 
        out[599] <= in[3293]; 
        out[600] <= in[2006]; 
        out[601] <= in[3693]; 
        out[602] <= in[3801]; 
        out[603] <= in[210]; 
        out[604] <= in[2877]; 
        out[605] <= in[3939]; 
        out[606] <= in[2784]; 
        out[607] <= in[3958]; 
        out[608] <= in[2271]; 
        out[609] <= in[1545]; 
        out[610] <= in[3153]; 
        out[611] <= in[815]; 
        out[612] <= in[1616]; 
        out[613] <= in[1122]; 
        out[614] <= in[721]; 
        out[615] <= in[133]; 
        out[616] <= in[3074]; 
        out[617] <= in[2959]; 
        out[618] <= in[1259]; 
        out[619] <= in[3339]; 
        out[620] <= in[86]; 
        out[621] <= in[2579]; 
        out[622] <= in[317]; 
        out[623] <= in[3696]; 
        out[624] <= in[2137]; 
        out[625] <= in[1330]; 
        out[626] <= in[1661]; 
        out[627] <= in[3039]; 
        out[628] <= in[123]; 
        out[629] <= in[2908]; 
        out[630] <= in[2290]; 
        out[631] <= in[1264]; 
        out[632] <= in[2652]; 
        out[633] <= in[1725]; 
        out[634] <= in[428]; 
        out[635] <= in[3150]; 
        out[636] <= in[3418]; 
        out[637] <= in[16]; 
        out[638] <= in[1760]; 
        out[639] <= in[3010]; 
        out[640] <= in[3264]; 
        out[641] <= in[3457]; 
        out[642] <= in[1176]; 
        out[643] <= in[2366]; 
        out[644] <= in[3234]; 
        out[645] <= in[2227]; 
        out[646] <= in[4036]; 
        out[647] <= in[425]; 
        out[648] <= in[3811]; 
        out[649] <= in[1929]; 
        out[650] <= in[879]; 
        out[651] <= in[1891]; 
        out[652] <= in[722]; 
        out[653] <= in[1492]; 
        out[654] <= in[1554]; 
        out[655] <= in[778]; 
        out[656] <= in[643]; 
        out[657] <= in[3185]; 
        out[658] <= in[3950]; 
        out[659] <= in[3143]; 
        out[660] <= in[526]; 
        out[661] <= in[177]; 
        out[662] <= in[1826]; 
        out[663] <= in[2632]; 
        out[664] <= in[2277]; 
        out[665] <= in[2311]; 
        out[666] <= in[358]; 
        out[667] <= in[1325]; 
        out[668] <= in[2558]; 
        out[669] <= in[877]; 
        out[670] <= in[1981]; 
        out[671] <= in[3079]; 
        out[672] <= in[2042]; 
        out[673] <= in[3902]; 
        out[674] <= in[1206]; 
        out[675] <= in[2256]; 
        out[676] <= in[941]; 
        out[677] <= in[1935]; 
        out[678] <= in[1513]; 
        out[679] <= in[1488]; 
        out[680] <= in[2437]; 
        out[681] <= in[3945]; 
        out[682] <= in[3372]; 
        out[683] <= in[1949]; 
        out[684] <= in[642]; 
        out[685] <= in[3403]; 
        out[686] <= in[1371]; 
        out[687] <= in[1612]; 
        out[688] <= in[1556]; 
        out[689] <= in[1188]; 
        out[690] <= in[700]; 
        out[691] <= in[3853]; 
        out[692] <= in[479]; 
        out[693] <= in[3218]; 
        out[694] <= in[518]; 
        out[695] <= in[1312]; 
        out[696] <= in[3084]; 
        out[697] <= in[1208]; 
        out[698] <= in[2340]; 
        out[699] <= in[3260]; 
        out[700] <= in[1261]; 
        out[701] <= in[2194]; 
        out[702] <= in[653]; 
        out[703] <= in[146]; 
        out[704] <= in[3179]; 
        out[705] <= in[2692]; 
        out[706] <= in[480]; 
        out[707] <= in[2036]; 
        out[708] <= in[187]; 
        out[709] <= in[3122]; 
        out[710] <= in[2800]; 
        out[711] <= in[937]; 
        out[712] <= in[3100]; 
        out[713] <= in[3189]; 
        out[714] <= in[2225]; 
        out[715] <= in[4037]; 
        out[716] <= in[998]; 
        out[717] <= in[460]; 
        out[718] <= in[3022]; 
        out[719] <= in[807]; 
        out[720] <= in[2677]; 
        out[721] <= in[508]; 
        out[722] <= in[1763]; 
        out[723] <= in[3050]; 
        out[724] <= in[2661]; 
        out[725] <= in[1012]; 
        out[726] <= in[69]; 
        out[727] <= in[1416]; 
        out[728] <= in[3743]; 
        out[729] <= in[1590]; 
        out[730] <= in[893]; 
        out[731] <= in[538]; 
        out[732] <= in[3427]; 
        out[733] <= in[694]; 
        out[734] <= in[789]; 
        out[735] <= in[3526]; 
        out[736] <= in[4052]; 
        out[737] <= in[3327]; 
        out[738] <= in[1960]; 
        out[739] <= in[2057]; 
        out[740] <= in[3399]; 
        out[741] <= in[3919]; 
        out[742] <= in[2099]; 
        out[743] <= in[2478]; 
        out[744] <= in[1921]; 
        out[745] <= in[2182]; 
        out[746] <= in[500]; 
        out[747] <= in[3701]; 
        out[748] <= in[1411]; 
        out[749] <= in[3322]; 
        out[750] <= in[3651]; 
        out[751] <= in[2471]; 
        out[752] <= in[3237]; 
        out[753] <= in[1924]; 
        out[754] <= in[2587]; 
        out[755] <= in[2030]; 
        out[756] <= in[4011]; 
        out[757] <= in[1712]; 
        out[758] <= in[206]; 
        out[759] <= in[714]; 
        out[760] <= in[1565]; 
        out[761] <= in[2739]; 
        out[762] <= in[1621]; 
        out[763] <= in[3586]; 
        out[764] <= in[53]; 
        out[765] <= in[2617]; 
        out[766] <= in[3424]; 
        out[767] <= in[968]; 
        out[768] <= in[523]; 
        out[769] <= in[3221]; 
        out[770] <= in[4035]; 
        out[771] <= in[2196]; 
        out[772] <= in[780]; 
        out[773] <= in[2731]; 
        out[774] <= in[3354]; 
        out[775] <= in[2508]; 
        out[776] <= in[3262]; 
        out[777] <= in[1022]; 
        out[778] <= in[2659]; 
        out[779] <= in[4079]; 
        out[780] <= in[3596]; 
        out[781] <= in[2672]; 
        out[782] <= in[3244]; 
        out[783] <= in[2777]; 
        out[784] <= in[3466]; 
        out[785] <= in[2916]; 
        out[786] <= in[3246]; 
        out[787] <= in[3289]; 
        out[788] <= in[1608]; 
        out[789] <= in[220]; 
        out[790] <= in[386]; 
        out[791] <= in[3898]; 
        out[792] <= in[1511]; 
        out[793] <= in[3135]; 
        out[794] <= in[599]; 
        out[795] <= in[1237]; 
        out[796] <= in[3456]; 
        out[797] <= in[357]; 
        out[798] <= in[4005]; 
        out[799] <= in[2090]; 
        out[800] <= in[108]; 
        out[801] <= in[630]; 
        out[802] <= in[408]; 
        out[803] <= in[2796]; 
        out[804] <= in[621]; 
        out[805] <= in[2874]; 
        out[806] <= in[531]; 
        out[807] <= in[2824]; 
        out[808] <= in[216]; 
        out[809] <= in[1385]; 
        out[810] <= in[2443]; 
        out[811] <= in[23]; 
        out[812] <= in[1815]; 
        out[813] <= in[7]; 
        out[814] <= in[2932]; 
        out[815] <= in[3700]; 
        out[816] <= in[1934]; 
        out[817] <= in[176]; 
        out[818] <= in[227]; 
        out[819] <= in[2174]; 
        out[820] <= in[1591]; 
        out[821] <= in[2436]; 
        out[822] <= in[1593]; 
        out[823] <= in[505]; 
        out[824] <= in[1380]; 
        out[825] <= in[4083]; 
        out[826] <= in[4041]; 
        out[827] <= in[2519]; 
        out[828] <= in[667]; 
        out[829] <= in[1887]; 
        out[830] <= in[4067]; 
        out[831] <= in[1690]; 
        out[832] <= in[3655]; 
        out[833] <= in[2403]; 
        out[834] <= in[1131]; 
        out[835] <= in[207]; 
        out[836] <= in[2027]; 
        out[837] <= in[3423]; 
        out[838] <= in[2274]; 
        out[839] <= in[63]; 
        out[840] <= in[2790]; 
        out[841] <= in[689]; 
        out[842] <= in[899]; 
        out[843] <= in[1870]; 
        out[844] <= in[3666]; 
        out[845] <= in[818]; 
        out[846] <= in[292]; 
        out[847] <= in[3782]; 
        out[848] <= in[84]; 
        out[849] <= in[3638]; 
        out[850] <= in[1539]; 
        out[851] <= in[2962]; 
        out[852] <= in[1460]; 
        out[853] <= in[1720]; 
        out[854] <= in[2656]; 
        out[855] <= in[461]; 
        out[856] <= in[2211]; 
        out[857] <= in[497]; 
        out[858] <= in[3692]; 
        out[859] <= in[314]; 
        out[860] <= in[1041]; 
        out[861] <= in[6]; 
        out[862] <= in[2917]; 
        out[863] <= in[3555]; 
        out[864] <= in[3281]; 
        out[865] <= in[2072]; 
        out[866] <= in[2514]; 
        out[867] <= in[1944]; 
        out[868] <= in[392]; 
        out[869] <= in[3518]; 
        out[870] <= in[1225]; 
        out[871] <= in[996]; 
        out[872] <= in[2146]; 
        out[873] <= in[4092]; 
        out[874] <= in[2260]; 
        out[875] <= in[1679]; 
        out[876] <= in[2681]; 
        out[877] <= in[3284]; 
        out[878] <= in[1027]; 
        out[879] <= in[959]; 
        out[880] <= in[3352]; 
        out[881] <= in[2577]; 
        out[882] <= in[3756]; 
        out[883] <= in[1696]; 
        out[884] <= in[138]; 
        out[885] <= in[1020]; 
        out[886] <= in[3467]; 
        out[887] <= in[786]; 
        out[888] <= in[2956]; 
        out[889] <= in[622]; 
        out[890] <= in[3587]; 
        out[891] <= in[3280]; 
        out[892] <= in[2402]; 
        out[893] <= in[3688]; 
        out[894] <= in[1977]; 
        out[895] <= in[3091]; 
        out[896] <= in[156]; 
        out[897] <= in[1464]; 
        out[898] <= in[2098]; 
        out[899] <= in[2658]; 
        out[900] <= in[634]; 
        out[901] <= in[0]; 
        out[902] <= in[862]; 
        out[903] <= in[347]; 
        out[904] <= in[349]; 
        out[905] <= in[1242]; 
        out[906] <= in[1836]; 
        out[907] <= in[1146]; 
        out[908] <= in[2832]; 
        out[909] <= in[636]; 
        out[910] <= in[535]; 
        out[911] <= in[3381]; 
        out[912] <= in[2535]; 
        out[913] <= in[475]; 
        out[914] <= in[3906]; 
        out[915] <= in[2791]; 
        out[916] <= in[2760]; 
        out[917] <= in[3432]; 
        out[918] <= in[2541]; 
        out[919] <= in[589]; 
        out[920] <= in[857]; 
        out[921] <= in[3834]; 
        out[922] <= in[1688]; 
        out[923] <= in[3663]; 
        out[924] <= in[2669]; 
        out[925] <= in[1903]; 
        out[926] <= in[115]; 
        out[927] <= in[1989]; 
        out[928] <= in[13]; 
        out[929] <= in[2387]; 
        out[930] <= in[1645]; 
        out[931] <= in[1456]; 
        out[932] <= in[1535]; 
        out[933] <= in[2899]; 
        out[934] <= in[1168]; 
        out[935] <= in[1494]; 
        out[936] <= in[4072]; 
        out[937] <= in[3337]; 
        out[938] <= in[1769]; 
        out[939] <= in[3239]; 
        out[940] <= in[3017]; 
        out[941] <= in[2772]; 
        out[942] <= in[1701]; 
        out[943] <= in[4031]; 
        out[944] <= in[294]; 
        out[945] <= in[1437]; 
        out[946] <= in[3859]; 
        out[947] <= in[983]; 
        out[948] <= in[1522]; 
        out[949] <= in[1641]; 
        out[950] <= in[3603]; 
        out[951] <= in[1523]; 
        out[952] <= in[2502]; 
        out[953] <= in[1192]; 
        out[954] <= in[2286]; 
        out[955] <= in[798]; 
        out[956] <= in[2152]; 
        out[957] <= in[253]; 
        out[958] <= in[1240]; 
        out[959] <= in[1118]; 
        out[960] <= in[3861]; 
        out[961] <= in[3935]; 
        out[962] <= in[2944]; 
        out[963] <= in[890]; 
        out[964] <= in[238]; 
        out[965] <= in[2805]; 
        out[966] <= in[3551]; 
        out[967] <= in[2590]; 
        out[968] <= in[905]; 
        out[969] <= in[3129]; 
        out[970] <= in[2678]; 
        out[971] <= in[644]; 
        out[972] <= in[3123]; 
        out[973] <= in[3021]; 
        out[974] <= in[2045]; 
        out[975] <= in[2255]; 
        out[976] <= in[1304]; 
        out[977] <= in[2037]; 
        out[978] <= in[2025]; 
        out[979] <= in[1987]; 
        out[980] <= in[3484]; 
        out[981] <= in[3335]; 
        out[982] <= in[1975]; 
        out[983] <= in[3407]; 
        out[984] <= in[1367]; 
        out[985] <= in[1638]; 
        out[986] <= in[3197]; 
        out[987] <= in[2534]; 
        out[988] <= in[791]; 
        out[989] <= in[3965]; 
        out[990] <= in[2516]; 
        out[991] <= in[2783]; 
        out[992] <= in[3080]; 
        out[993] <= in[898]; 
        out[994] <= in[277]; 
        out[995] <= in[2201]; 
        out[996] <= in[1917]; 
        out[997] <= in[3607]; 
        out[998] <= in[955]; 
        out[999] <= in[1401]; 
        out[1000] <= in[874]; 
        out[1001] <= in[2422]; 
        out[1002] <= in[437]; 
        out[1003] <= in[3496]; 
        out[1004] <= in[614]; 
        out[1005] <= in[2082]; 
        out[1006] <= in[1843]; 
        out[1007] <= in[2640]; 
        out[1008] <= in[3675]; 
        out[1009] <= in[3671]; 
        out[1010] <= in[36]; 
        out[1011] <= in[3884]; 
        out[1012] <= in[217]; 
        out[1013] <= in[1749]; 
        out[1014] <= in[2315]; 
        out[1015] <= in[1229]; 
        out[1016] <= in[3490]; 
        out[1017] <= in[2209]; 
        out[1018] <= in[1021]; 
        out[1019] <= in[2744]; 
        out[1020] <= in[368]; 
        out[1021] <= in[972]; 
        out[1022] <= in[534]; 
        out[1023] <= in[2475]; 
        out[1024] <= in[3744]; 
        out[1025] <= in[3924]; 
        out[1026] <= in[3765]; 
        out[1027] <= in[3625]; 
        out[1028] <= in[1289]; 
        out[1029] <= in[1448]; 
        out[1030] <= in[2113]; 
        out[1031] <= in[2477]; 
        out[1032] <= in[3595]; 
        out[1033] <= in[1440]; 
        out[1034] <= in[1317]; 
        out[1035] <= in[3548]; 
        out[1036] <= in[3639]; 
        out[1037] <= in[1472]; 
        out[1038] <= in[978]; 
        out[1039] <= in[2513]; 
        out[1040] <= in[2018]; 
        out[1041] <= in[943]; 
        out[1042] <= in[8]; 
        out[1043] <= in[1247]; 
        out[1044] <= in[3308]; 
        out[1045] <= in[3498]; 
        out[1046] <= in[162]; 
        out[1047] <= in[3857]; 
        out[1048] <= in[840]; 
        out[1049] <= in[2573]; 
        out[1050] <= in[631]; 
        out[1051] <= in[3827]; 
        out[1052] <= in[1110]; 
        out[1053] <= in[2032]; 
        out[1054] <= in[1275]; 
        out[1055] <= in[3515]; 
        out[1056] <= in[3229]; 
        out[1057] <= in[2061]; 
        out[1058] <= in[1717]; 
        out[1059] <= in[14]; 
        out[1060] <= in[2183]; 
        out[1061] <= in[3047]; 
        out[1062] <= in[3993]; 
        out[1063] <= in[376]; 
        out[1064] <= in[3728]; 
        out[1065] <= in[2005]; 
        out[1066] <= in[3401]; 
        out[1067] <= in[2050]; 
        out[1068] <= in[3917]; 
        out[1069] <= in[2088]; 
        out[1070] <= in[3358]; 
        out[1071] <= in[2952]; 
        out[1072] <= in[3778]; 
        out[1073] <= in[254]; 
        out[1074] <= in[3031]; 
        out[1075] <= in[1175]; 
        out[1076] <= in[192]; 
        out[1077] <= in[1326]; 
        out[1078] <= in[444]; 
        out[1079] <= in[2935]; 
        out[1080] <= in[450]; 
        out[1081] <= in[285]; 
        out[1082] <= in[3194]; 
        out[1083] <= in[1907]; 
        out[1084] <= in[2770]; 
        out[1085] <= in[1489]; 
        out[1086] <= in[12]; 
        out[1087] <= in[1438]; 
        out[1088] <= in[596]; 
        out[1089] <= in[716]; 
        out[1090] <= in[963]; 
        out[1091] <= in[3077]; 
        out[1092] <= in[2221]; 
        out[1093] <= in[2829]; 
        out[1094] <= in[3646]; 
        out[1095] <= in[2693]; 
        out[1096] <= in[35]; 
        out[1097] <= in[2193]; 
        out[1098] <= in[880]; 
        out[1099] <= in[2754]; 
        out[1100] <= in[1496]; 
        out[1101] <= in[687]; 
        out[1102] <= in[3583]; 
        out[1103] <= in[3094]; 
        out[1104] <= in[1282]; 
        out[1105] <= in[2643]; 
        out[1106] <= in[1615]; 
        out[1107] <= in[3912]; 
        out[1108] <= in[1569]; 
        out[1109] <= in[749]; 
        out[1110] <= in[3726]; 
        out[1111] <= in[1541]; 
        out[1112] <= in[2188]; 
        out[1113] <= in[3864]; 
        out[1114] <= in[524]; 
        out[1115] <= in[3867]; 
        out[1116] <= in[3716]; 
        out[1117] <= in[673]; 
        out[1118] <= in[3809]; 
        out[1119] <= in[2909]; 
        out[1120] <= in[3571]; 
        out[1121] <= in[3062]; 
        out[1122] <= in[2457]; 
        out[1123] <= in[2680]; 
        out[1124] <= in[3087]; 
        out[1125] <= in[2776]; 
        out[1126] <= in[82]; 
        out[1127] <= in[914]; 
        out[1128] <= in[4091]; 
        out[1129] <= in[1249]; 
        out[1130] <= in[1718]; 
        out[1131] <= in[3627]; 
        out[1132] <= in[3979]; 
        out[1133] <= in[3943]; 
        out[1134] <= in[3111]; 
        out[1135] <= in[1898]; 
        out[1136] <= in[1001]; 
        out[1137] <= in[2368]; 
        out[1138] <= in[173]; 
        out[1139] <= in[897]; 
        out[1140] <= in[3529]; 
        out[1141] <= in[4048]; 
        out[1142] <= in[2548]; 
        out[1143] <= in[2743]; 
        out[1144] <= in[313]; 
        out[1145] <= in[157]; 
        out[1146] <= in[1290]; 
        out[1147] <= in[2058]; 
        out[1148] <= in[198]; 
        out[1149] <= in[200]; 
        out[1150] <= in[575]; 
        out[1151] <= in[2011]; 
        out[1152] <= in[1603]; 
        out[1153] <= in[2285]; 
        out[1154] <= in[1184]; 
        out[1155] <= in[1682]; 
        out[1156] <= in[1430]; 
        out[1157] <= in[806]; 
        out[1158] <= in[763]; 
        out[1159] <= in[1684]; 
        out[1160] <= in[1952]; 
        out[1161] <= in[2876]; 
        out[1162] <= in[734]; 
        out[1163] <= in[3222]; 
        out[1164] <= in[4085]; 
        out[1165] <= in[3597]; 
        out[1166] <= in[2825]; 
        out[1167] <= in[112]; 
        out[1168] <= in[2016]; 
        out[1169] <= in[2360]; 
        out[1170] <= in[2008]; 
        out[1171] <= in[3092]; 
        out[1172] <= in[3883]; 
        out[1173] <= in[4073]; 
        out[1174] <= in[3925]; 
        out[1175] <= in[2851]; 
        out[1176] <= in[1505]; 
        out[1177] <= in[3506]; 
        out[1178] <= in[3545]; 
        out[1179] <= in[2627]; 
        out[1180] <= in[1144]; 
        out[1181] <= in[1649]; 
        out[1182] <= in[852]; 
        out[1183] <= in[1681]; 
        out[1184] <= in[4062]; 
        out[1185] <= in[4014]; 
        out[1186] <= in[2109]; 
        out[1187] <= in[3063]; 
        out[1188] <= in[1715]; 
        out[1189] <= in[892]; 
        out[1190] <= in[1062]; 
        out[1191] <= in[3317]; 
        out[1192] <= in[1273]; 
        out[1193] <= in[1534]; 
        out[1194] <= in[974]; 
        out[1195] <= in[3453]; 
        out[1196] <= in[4042]; 
        out[1197] <= in[1026]; 
        out[1198] <= in[675]; 
        out[1199] <= in[2814]; 
        out[1200] <= in[3605]; 
        out[1201] <= in[565]; 
        out[1202] <= in[2826]; 
        out[1203] <= in[863]; 
        out[1204] <= in[602]; 
        out[1205] <= in[704]; 
        out[1206] <= in[1867]; 
        out[1207] <= in[3376]; 
        out[1208] <= in[111]; 
        out[1209] <= in[3579]; 
        out[1210] <= in[826]; 
        out[1211] <= in[1838]; 
        out[1212] <= in[3342]; 
        out[1213] <= in[1572]; 
        out[1214] <= in[1166]; 
        out[1215] <= in[3018]; 
        out[1216] <= in[607]; 
        out[1217] <= in[1651]; 
        out[1218] <= in[3422]; 
        out[1219] <= in[2622]; 
        out[1220] <= in[312]; 
        out[1221] <= in[2871]; 
        out[1222] <= in[3097]; 
        out[1223] <= in[3076]; 
        out[1224] <= in[2363]; 
        out[1225] <= in[1126]; 
        out[1226] <= in[1776]; 
        out[1227] <= in[3951]; 
        out[1228] <= in[297]; 
        out[1229] <= in[2461]; 
        out[1230] <= in[3561]; 
        out[1231] <= in[770]; 
        out[1232] <= in[3235]; 
        out[1233] <= in[3888]; 
        out[1234] <= in[1816]; 
        out[1235] <= in[2882]; 
        out[1236] <= in[1819]; 
        out[1237] <= in[2215]; 
        out[1238] <= in[3029]; 
        out[1239] <= in[3916]; 
        out[1240] <= in[3203]; 
        out[1241] <= in[2690]; 
        out[1242] <= in[3871]; 
        out[1243] <= in[418]; 
        out[1244] <= in[2687]; 
        out[1245] <= in[554]; 
        out[1246] <= in[3042]; 
        out[1247] <= in[1382]; 
        out[1248] <= in[340]; 
        out[1249] <= in[2170]; 
        out[1250] <= in[178]; 
        out[1251] <= in[440]; 
        out[1252] <= in[1220]; 
        out[1253] <= in[1965]; 
        out[1254] <= in[3251]; 
        out[1255] <= in[3880]; 
        out[1256] <= in[2416]; 
        out[1257] <= in[1136]; 
        out[1258] <= in[1163]; 
        out[1259] <= in[2308]; 
        out[1260] <= in[2305]; 
        out[1261] <= in[3175]; 
        out[1262] <= in[2230]; 
        out[1263] <= in[1156]; 
        out[1264] <= in[3821]; 
        out[1265] <= in[2976]; 
        out[1266] <= in[288]; 
        out[1267] <= in[1553]; 
        out[1268] <= in[1791]; 
        out[1269] <= in[1000]; 
        out[1270] <= in[2167]; 
        out[1271] <= in[1667]; 
        out[1272] <= in[2143]; 
        out[1273] <= in[124]; 
        out[1274] <= in[2357]; 
        out[1275] <= in[1963]; 
        out[1276] <= in[3723]; 
        out[1277] <= in[2531]; 
        out[1278] <= in[1170]; 
        out[1279] <= in[3083]; 
        out[1280] <= in[3386]; 
        out[1281] <= in[1093]; 
        out[1282] <= in[2848]; 
        out[1283] <= in[3355]; 
        out[1284] <= in[2122]; 
        out[1285] <= in[856]; 
        out[1286] <= in[1316]; 
        out[1287] <= in[2948]; 
        out[1288] <= in[3305]; 
        out[1289] <= in[2540]; 
        out[1290] <= in[2887]; 
        out[1291] <= in[3885]; 
        out[1292] <= in[3628]; 
        out[1293] <= in[4045]; 
        out[1294] <= in[1959]; 
        out[1295] <= in[2200]; 
        out[1296] <= in[75]; 
        out[1297] <= in[1265]; 
        out[1298] <= in[2118]; 
        out[1299] <= in[1829]; 
        out[1300] <= in[1375]; 
        out[1301] <= in[4017]; 
        out[1302] <= in[829]; 
        out[1303] <= in[401]; 
        out[1304] <= in[1069]; 
        out[1305] <= in[953]; 
        out[1306] <= in[360]; 
        out[1307] <= in[2942]; 
        out[1308] <= in[3370]; 
        out[1309] <= in[3028]; 
        out[1310] <= in[2392]; 
        out[1311] <= in[2999]; 
        out[1312] <= in[956]; 
        out[1313] <= in[1630]; 
        out[1314] <= in[1415]; 
        out[1315] <= in[2737]; 
        out[1316] <= in[743]; 
        out[1317] <= in[4012]; 
        out[1318] <= in[572]; 
        out[1319] <= in[1610]; 
        out[1320] <= in[584]; 
        out[1321] <= in[717]; 
        out[1322] <= in[2244]; 
        out[1323] <= in[2978]; 
        out[1324] <= in[3415]; 
        out[1325] <= in[1221]; 
        out[1326] <= in[2080]; 
        out[1327] <= in[2401]; 
        out[1328] <= in[1169]; 
        out[1329] <= in[3787]; 
        out[1330] <= in[3720]; 
        out[1331] <= in[296]; 
        out[1332] <= in[1368]; 
        out[1333] <= in[2756]; 
        out[1334] <= in[3148]; 
        out[1335] <= in[1467]; 
        out[1336] <= in[3009]; 
        out[1337] <= in[2705]; 
        out[1338] <= in[946]; 
        out[1339] <= in[2377]; 
        out[1340] <= in[3273]; 
        out[1341] <= in[907]; 
        out[1342] <= in[2365]; 
        out[1343] <= in[1779]; 
        out[1344] <= in[366]; 
        out[1345] <= in[1711]; 
        out[1346] <= in[3272]; 
        out[1347] <= in[2895]; 
        out[1348] <= in[2889]; 
        out[1349] <= in[2504]; 
        out[1350] <= in[648]; 
        out[1351] <= in[1253]; 
        out[1352] <= in[502]; 
        out[1353] <= in[3236]; 
        out[1354] <= in[1994]; 
        out[1355] <= in[2581]; 
        out[1356] <= in[3522]; 
        out[1357] <= in[615]; 
        out[1358] <= in[1199]; 
        out[1359] <= in[958]; 
        out[1360] <= in[68]; 
        out[1361] <= in[1660]; 
        out[1362] <= in[2103]; 
        out[1363] <= in[130]; 
        out[1364] <= in[3184]; 
        out[1365] <= in[2779]; 
        out[1366] <= in[1268]; 
        out[1367] <= in[3602]; 
        out[1368] <= in[2552]; 
        out[1369] <= in[1999]; 
        out[1370] <= in[1894]; 
        out[1371] <= in[1915]; 
        out[1372] <= in[659]; 
        out[1373] <= in[4027]; 
        out[1374] <= in[1753]; 
        out[1375] <= in[1498]; 
        out[1376] <= in[2961]; 
        out[1377] <= in[2280]; 
        out[1378] <= in[2566]; 
        out[1379] <= in[3788]; 
        out[1380] <= in[679]; 
        out[1381] <= in[3686]; 
        out[1382] <= in[397]; 
        out[1383] <= in[3685]; 
        out[1384] <= in[3577]; 
        out[1385] <= in[2641]; 
        out[1386] <= in[1939]; 
        out[1387] <= in[3449]; 
        out[1388] <= in[1525]; 
        out[1389] <= in[1413]; 
        out[1390] <= in[865]; 
        out[1391] <= in[1914]; 
        out[1392] <= in[213]; 
        out[1393] <= in[748]; 
        out[1394] <= in[331]; 
        out[1395] <= in[906]; 
        out[1396] <= in[1086]; 
        out[1397] <= in[3580]; 
        out[1398] <= in[421]; 
        out[1399] <= in[2919]; 
        out[1400] <= in[3434]; 
        out[1401] <= in[3921]; 
        out[1402] <= in[3149]; 
        out[1403] <= in[2329]; 
        out[1404] <= in[143]; 
        out[1405] <= in[1532]; 
        out[1406] <= in[3016]; 
        out[1407] <= in[3703]; 
        out[1408] <= in[878]; 
        out[1409] <= in[1284]; 
        out[1410] <= in[99]; 
        out[1411] <= in[3661]; 
        out[1412] <= in[1376]; 
        out[1413] <= in[4022]; 
        out[1414] <= in[3904]; 
        out[1415] <= in[1751]; 
        out[1416] <= in[1286]; 
        out[1417] <= in[1662]; 
        out[1418] <= in[85]; 
        out[1419] <= in[352]; 
        out[1420] <= in[3737]; 
        out[1421] <= in[986]; 
        out[1422] <= in[2884]; 
        out[1423] <= in[183]; 
        out[1424] <= in[1255]; 
        out[1425] <= in[438]; 
        out[1426] <= in[3707]; 
        out[1427] <= in[184]; 
        out[1428] <= in[3584]; 
        out[1429] <= in[1479]; 
        out[1430] <= in[1137]; 
        out[1431] <= in[3187]; 
        out[1432] <= in[541]; 
        out[1433] <= in[2013]; 
        out[1434] <= in[2822]; 
        out[1435] <= in[603]; 
        out[1436] <= in[649]; 
        out[1437] <= in[723]; 
        out[1438] <= in[1521]; 
        out[1439] <= in[3795]; 
        out[1440] <= in[2898]; 
        out[1441] <= in[1426]; 
        out[1442] <= in[3053]; 
        out[1443] <= in[2755]; 
        out[1444] <= in[2860]; 
        out[1445] <= in[2616]; 
        out[1446] <= in[3307]; 
        out[1447] <= in[1015]; 
        out[1448] <= in[2409]; 
        out[1449] <= in[94]; 
        out[1450] <= in[2650]; 
        out[1451] <= in[2460]; 
        out[1452] <= in[48]; 
        out[1453] <= in[761]; 
        out[1454] <= in[131]; 
        out[1455] <= in[2145]; 
        out[1456] <= in[306]; 
        out[1457] <= in[3011]; 
        out[1458] <= in[612]; 
        out[1459] <= in[3452]; 
        out[1460] <= in[459]; 
        out[1461] <= in[3835]; 
        out[1462] <= in[1731]; 
        out[1463] <= in[2456]; 
        out[1464] <= in[299]; 
        out[1465] <= in[1582]; 
        out[1466] <= in[1336]; 
        out[1467] <= in[193]; 
        out[1468] <= in[510]; 
        out[1469] <= in[134]; 
        out[1470] <= in[3020]; 
        out[1471] <= in[812]; 
        out[1472] <= in[2761]; 
        out[1473] <= in[1353]; 
        out[1474] <= in[3761]; 
        out[1475] <= in[3826]; 
        out[1476] <= in[1970]; 
        out[1477] <= in[3822]; 
        out[1478] <= in[1571]; 
        out[1479] <= in[973]; 
        out[1480] <= in[1044]; 
        out[1481] <= in[3114]; 
        out[1482] <= in[3878]; 
        out[1483] <= in[3574]; 
        out[1484] <= in[3183]; 
        out[1485] <= in[4050]; 
        out[1486] <= in[2446]; 
        out[1487] <= in[2647]; 
        out[1488] <= in[2476]; 
        out[1489] <= in[3267]; 
        out[1490] <= in[1575]; 
        out[1491] <= in[3363]; 
        out[1492] <= in[708]; 
        out[1493] <= in[1030]; 
        out[1494] <= in[1150]; 
        out[1495] <= in[1938]; 
        out[1496] <= in[231]; 
        out[1497] <= in[2964]; 
        out[1498] <= in[149]; 
        out[1499] <= in[2571]; 
        out[1500] <= in[417]; 
        out[1501] <= in[1544]; 
        out[1502] <= in[410]; 
        out[1503] <= in[2131]; 
        out[1504] <= in[4053]; 
        out[1505] <= in[3717]; 
        out[1506] <= in[1750]; 
        out[1507] <= in[674]; 
        out[1508] <= in[2139]; 
        out[1509] <= in[758]; 
        out[1510] <= in[3739]; 
        out[1511] <= in[1332]; 
        out[1512] <= in[2325]; 
        out[1513] <= in[3003]; 
        out[1514] <= in[1471]; 
        out[1515] <= in[2073]; 
        out[1516] <= in[516]; 
        out[1517] <= in[4002]; 
        out[1518] <= in[1920]; 
        out[1519] <= in[1798]; 
        out[1520] <= in[281]; 
        out[1521] <= in[1238]; 
        out[1522] <= in[3421]; 
        out[1523] <= in[2715]; 
        out[1524] <= in[1509]; 
        out[1525] <= in[831]; 
        out[1526] <= in[2473]; 
        out[1527] <= in[2890]; 
        out[1528] <= in[662]; 
        out[1529] <= in[2536]; 
        out[1530] <= in[1730]; 
        out[1531] <= in[1370]; 
        out[1532] <= in[3347]; 
        out[1533] <= in[3410]; 
        out[1534] <= in[585]; 
        out[1535] <= in[3443]; 
        out[1536] <= in[557]; 
        out[1537] <= in[1800]; 
        out[1538] <= in[343]; 
        out[1539] <= in[3055]; 
        out[1540] <= in[3380]; 
        out[1541] <= in[321]; 
        out[1542] <= in[1239]; 
        out[1543] <= in[3590]; 
        out[1544] <= in[1420]; 
        out[1545] <= in[2843]; 
        out[1546] <= in[1484]; 
        out[1547] <= in[2081]; 
        out[1548] <= in[1281]; 
        out[1549] <= in[3182]; 
        out[1550] <= in[350]; 
        out[1551] <= in[1315]; 
        out[1552] <= in[837]; 
        out[1553] <= in[1292]; 
        out[1554] <= in[2171]; 
        out[1555] <= in[2979]; 
        out[1556] <= in[379]; 
        out[1557] <= in[458]; 
        out[1558] <= in[3931]; 
        out[1559] <= in[1014]; 
        out[1560] <= in[771]; 
        out[1561] <= in[2054]; 
        out[1562] <= in[3471]; 
        out[1563] <= in[1883]; 
        out[1564] <= in[1605]; 
        out[1565] <= in[3558]; 
        out[1566] <= in[3278]; 
        out[1567] <= in[3976]; 
        out[1568] <= in[1073]; 
        out[1569] <= in[1581]; 
        out[1570] <= in[3961]; 
        out[1571] <= in[3905]; 
        out[1572] <= in[2239]; 
        out[1573] <= in[1222]; 
        out[1574] <= in[426]; 
        out[1575] <= in[1595]; 
        out[1576] <= in[2275]; 
        out[1577] <= in[58]; 
        out[1578] <= in[3749]; 
        out[1579] <= in[949]; 
        out[1580] <= in[2218]; 
        out[1581] <= in[2934]; 
        out[1582] <= in[64]; 
        out[1583] <= in[3261]; 
        out[1584] <= in[3733]; 
        out[1585] <= in[3425]; 
        out[1586] <= in[3706]; 
        out[1587] <= in[1394]; 
        out[1588] <= in[439]; 
        out[1589] <= in[4063]; 
        out[1590] <= in[1895]; 
        out[1591] <= in[1451]; 
        out[1592] <= in[3446]; 
        out[1593] <= in[1627]; 
        out[1594] <= in[362]; 
        out[1595] <= in[1656]; 
        out[1596] <= in[2811]; 
        out[1597] <= in[2427]; 
        out[1598] <= in[3539]; 
        out[1599] <= in[1010]; 
        out[1600] <= in[2938]; 
        out[1601] <= in[2163]; 
        out[1602] <= in[405]; 
        out[1603] <= in[3318]; 
        out[1604] <= in[4049]; 
        out[1605] <= in[2208]; 
        out[1606] <= in[2370]; 
        out[1607] <= in[481]; 
        out[1608] <= in[3458]; 
        out[1609] <= in[87]; 
        out[1610] <= in[2563]; 
        out[1611] <= in[476]; 
        out[1612] <= in[3275]; 
        out[1613] <= in[2059]; 
        out[1614] <= in[1613]; 
        out[1615] <= in[1051]; 
        out[1616] <= in[2608]; 
        out[1617] <= in[1568]; 
        out[1618] <= in[3644]; 
        out[1619] <= in[1884]; 
        out[1620] <= in[3059]; 
        out[1621] <= in[4068]; 
        out[1622] <= in[2445]; 
        out[1623] <= in[4060]; 
        out[1624] <= in[3450]; 
        out[1625] <= in[2667]; 
        out[1626] <= in[3901]; 
        out[1627] <= in[1853]; 
        out[1628] <= in[2389]; 
        out[1629] <= in[1787]; 
        out[1630] <= in[179]; 
        out[1631] <= in[2134]; 
        out[1632] <= in[251]; 
        out[1633] <= in[3704]; 
        out[1634] <= in[809]; 
        out[1635] <= in[836]; 
        out[1636] <= in[917]; 
        out[1637] <= in[2542]; 
        out[1638] <= in[2198]; 
        out[1639] <= in[2270]; 
        out[1640] <= in[2856]; 
        out[1641] <= in[1490]; 
        out[1642] <= in[2108]; 
        out[1643] <= in[1466]; 
        out[1644] <= in[150]; 
        out[1645] <= in[2518]; 
        out[1646] <= in[2599]; 
        out[1647] <= in[847]; 
        out[1648] <= in[2254]; 
        out[1649] <= in[651]; 
        out[1650] <= in[2747]; 
        out[1651] <= in[3340]; 
        out[1652] <= in[2390]; 
        out[1653] <= in[3286]; 
        out[1654] <= in[2888]; 
        out[1655] <= in[214]; 
        out[1656] <= in[2698]; 
        out[1657] <= in[868]; 
        out[1658] <= in[1721]; 
        out[1659] <= in[336]; 
        out[1660] <= in[855]; 
        out[1661] <= in[2655]; 
        out[1662] <= in[1]; 
        out[1663] <= in[323]; 
        out[1664] <= in[2937]; 
        out[1665] <= in[2490]; 
        out[1666] <= in[2128]; 
        out[1667] <= in[393]; 
        out[1668] <= in[3566]; 
        out[1669] <= in[3687]; 
        out[1670] <= in[1879]; 
        out[1671] <= in[10]; 
        out[1672] <= in[1697]; 
        out[1673] <= in[3755]; 
        out[1674] <= in[1566]; 
        out[1675] <= in[773]; 
        out[1676] <= in[245]; 
        out[1677] <= in[1973]; 
        out[1678] <= in[2375]; 
        out[1679] <= in[1743]; 
        out[1680] <= in[2240]; 
        out[1681] <= in[1162]; 
        out[1682] <= in[259]; 
        out[1683] <= in[2723]; 
        out[1684] <= in[436]; 
        out[1685] <= in[577]; 
        out[1686] <= in[3698]; 
        out[1687] <= in[2079]; 
        out[1688] <= in[2880]; 
        out[1689] <= in[1871]; 
        out[1690] <= in[797]; 
        out[1691] <= in[2921]; 
        out[1692] <= in[3497]; 
        out[1693] <= in[234]; 
        out[1694] <= in[895]; 
        out[1695] <= in[3023]; 
        out[1696] <= in[1536]; 
        out[1697] <= in[3125]; 
        out[1698] <= in[1195]; 
        out[1699] <= in[3672]; 
        out[1700] <= in[258]; 
        out[1701] <= in[303]; 
        out[1702] <= in[792]; 
        out[1703] <= in[1034]; 
        out[1704] <= in[4087]; 
        out[1705] <= in[2318]; 
        out[1706] <= in[618]; 
        out[1707] <= in[1243]; 
        out[1708] <= in[2266]; 
        out[1709] <= in[3404]; 
        out[1710] <= in[1311]; 
        out[1711] <= in[591]; 
        out[1712] <= in[2249]; 
        out[1713] <= in[3576]; 
        out[1714] <= in[3572]; 
        out[1715] <= in[3632]; 
        out[1716] <= in[2284]; 
        out[1717] <= in[101]; 
        out[1718] <= in[2828]; 
        out[1719] <= in[211]; 
        out[1720] <= in[2019]; 
        out[1721] <= in[1210]; 
        out[1722] <= in[3819]; 
        out[1723] <= in[3048]; 
        out[1724] <= in[3109]; 
        out[1725] <= in[1056]; 
        out[1726] <= in[3892]; 
        out[1727] <= in[1061]; 
        out[1728] <= in[228]; 
        out[1729] <= in[3792]; 
        out[1730] <= in[2553]; 
        out[1731] <= in[711]; 
        out[1732] <= in[3684]; 
        out[1733] <= in[3598]; 
        out[1734] <= in[1586]; 
        out[1735] <= in[1765]; 
        out[1736] <= in[1307]; 
        out[1737] <= in[3015]; 
        out[1738] <= in[2205]; 
        out[1739] <= in[598]; 
        out[1740] <= in[2559]; 
        out[1741] <= in[1832]; 
        out[1742] <= in[2901]; 
        out[1743] <= in[4]; 
        out[1744] <= in[3377]; 
        out[1745] <= in[1497]; 
        out[1746] <= in[3108]; 
        out[1747] <= in[1607]; 
        out[1748] <= in[2855]; 
        out[1749] <= in[3492]; 
        out[1750] <= in[581]; 
        out[1751] <= in[698]; 
        out[1752] <= in[537]; 
        out[1753] <= in[2430]; 
        out[1754] <= in[2074]; 
        out[1755] <= in[2164]; 
        out[1756] <= in[3604]; 
        out[1757] <= in[2452]; 
        out[1758] <= in[3113]; 
        out[1759] <= in[3903]; 
        out[1760] <= in[1418]; 
        out[1761] <= in[2555]; 
        out[1762] <= in[1224]; 
        out[1763] <= in[2233]; 
        out[1764] <= in[3412]; 
        out[1765] <= in[2424]; 
        out[1766] <= in[1654]; 
        out[1767] <= in[1419]; 
        out[1768] <= in[2292]; 
        out[1769] <= in[104]; 
        out[1770] <= in[3255]; 
        out[1771] <= in[2455]; 
        out[1772] <= in[2077]; 
        out[1773] <= in[2545]; 
        out[1774] <= in[889]; 
        out[1775] <= in[1378]; 
        out[1776] <= in[2787]; 
        out[1777] <= in[1606]; 
        out[1778] <= in[660]; 
        out[1779] <= in[4018]; 
        out[1780] <= in[141]; 
        out[1781] <= in[620]; 
        out[1782] <= in[424]; 
        out[1783] <= in[3856]; 
        out[1784] <= in[1642]; 
        out[1785] <= in[32]; 
        out[1786] <= in[4007]; 
        out[1787] <= in[962]; 
        out[1788] <= in[1587]; 
        out[1789] <= in[3201]; 
        out[1790] <= in[3523]; 
        out[1791] <= in[2380]; 
        out[1792] <= in[2689]; 
        out[1793] <= in[736]; 
        out[1794] <= in[2636]; 
        out[1795] <= in[3205]; 
        out[1796] <= in[2421]; 
        out[1797] <= in[816]; 
        out[1798] <= in[3828]; 
        out[1799] <= in[1704]; 
        out[1800] <= in[3369]; 
        out[1801] <= in[1781]; 
        out[1802] <= in[3913]; 
        out[1803] <= in[11]; 
        out[1804] <= in[1992]; 
        out[1805] <= in[1331]; 
        out[1806] <= in[3968]; 
        out[1807] <= in[2301]; 
        out[1808] <= in[3527]; 
        out[1809] <= in[737]; 
        out[1810] <= in[1159]; 
        out[1811] <= in[97]; 
        out[1812] <= in[3411]; 
        out[1813] <= in[2592]; 
        out[1814] <= in[3673]; 
        out[1815] <= in[586]; 
        out[1816] <= in[808]; 
        out[1817] <= in[1480]; 
        out[1818] <= in[166]; 
        out[1819] <= in[3800]; 
        out[1820] <= in[100]; 
        out[1821] <= in[4095]; 
        out[1822] <= in[399]; 
        out[1823] <= in[715]; 
        out[1824] <= in[327]; 
        out[1825] <= in[1075]; 
        out[1826] <= in[2896]; 
        out[1827] <= in[3438]; 
        out[1828] <= in[1308]; 
        out[1829] <= in[1962]; 
        out[1830] <= in[1241]; 
        out[1831] <= in[1623]; 
        out[1832] <= in[1343]; 
        out[1833] <= in[709]; 
        out[1834] <= in[2353]; 
        out[1835] <= in[4082]; 
        out[1836] <= in[3294]; 
        out[1837] <= in[875]; 
        out[1838] <= in[1257]; 
        out[1839] <= in[606]; 
        out[1840] <= in[1945]; 
        out[1841] <= in[2406]; 
        out[1842] <= in[819]; 
        out[1843] <= in[223]; 
        out[1844] <= in[443]; 
        out[1845] <= in[3190]; 
        out[1846] <= in[2206]; 
        out[1847] <= in[1722]; 
        out[1848] <= in[858]; 
        out[1849] <= in[1888]; 
        out[1850] <= in[2313]; 
        out[1851] <= in[3689]; 
        out[1852] <= in[3338]; 
        out[1853] <= in[1771]; 
        out[1854] <= in[1872]; 
        out[1855] <= in[1812]; 
        out[1856] <= in[720]; 
        out[1857] <= in[3563]; 
        out[1858] <= in[2087]; 
        out[1859] <= in[3842]; 
        out[1860] <= in[632]; 
        out[1861] <= in[1777]; 
        out[1862] <= in[2930]; 
        out[1863] <= in[2736]; 
        out[1864] <= in[628]; 
        out[1865] <= in[121]; 
        out[1866] <= in[601]; 
        out[1867] <= in[3932]; 
        out[1868] <= in[1454]; 
        out[1869] <= in[564]; 
        out[1870] <= in[4008]; 
        out[1871] <= in[583]; 
        out[1872] <= in[2369]; 
        out[1873] <= in[965]; 
        out[1874] <= in[665]; 
        out[1875] <= in[2135]; 
        out[1876] <= in[433]; 
        out[1877] <= in[2820]; 
        out[1878] <= in[3374]; 
        out[1879] <= in[1567]; 
        out[1880] <= in[2966]; 
        out[1881] <= in[3978]; 
        out[1882] <= in[3564]; 
        out[1883] <= in[2014]; 
        out[1884] <= in[2328]; 
        out[1885] <= in[1911]; 
        out[1886] <= in[1547]; 
        out[1887] <= in[3784]; 
        out[1888] <= in[3775]; 
        out[1889] <= in[181]; 
        out[1890] <= in[1848]; 
        out[1891] <= in[1452]; 
        out[1892] <= in[1417]; 
        out[1893] <= in[2120]; 
        out[1894] <= in[310]; 
        out[1895] <= in[1529]; 
        out[1896] <= in[2383]; 
        out[1897] <= in[1059]; 
        out[1898] <= in[3008]; 
        out[1899] <= in[2147]; 
        out[1900] <= in[345]; 
        out[1901] <= in[2806]; 
        out[1902] <= in[2133]; 
        out[1903] <= in[2530]; 
        out[1904] <= in[827]; 
        out[1905] <= in[273]; 
        out[1906] <= in[3214]; 
        out[1907] <= in[1925]; 
        out[1908] <= in[1406]; 
        out[1909] <= in[169]; 
        out[1910] <= in[1528]; 
        out[1911] <= in[3191]; 
        out[1912] <= in[3808]; 
        out[1913] <= in[1735]; 
        out[1914] <= in[28]; 
        out[1915] <= in[391]; 
        out[1916] <= in[190]; 
        out[1917] <= in[2773]; 
        out[1918] <= in[2498]; 
        out[1919] <= in[1830]; 
        out[1920] <= in[2686]; 
        out[1921] <= in[4059]; 
        out[1922] <= in[1178]; 
        out[1923] <= in[2853]; 
        out[1924] <= in[2586]; 
        out[1925] <= in[677]; 
        out[1926] <= in[269]; 
        out[1927] <= in[2489]; 
        out[1928] <= in[148]; 
        out[1929] <= in[1102]; 
        out[1930] <= in[491]; 
        out[1931] <= in[1119]; 
        out[1932] <= in[1618]; 
        out[1933] <= in[776]; 
        out[1934] <= in[2356]; 
        out[1935] <= in[224]; 
        out[1936] <= in[490]; 
        out[1937] <= in[511]; 
        out[1938] <= in[886]; 
        out[1939] <= in[1979]; 
        out[1940] <= in[2217]; 
        out[1941] <= in[2838]; 
        out[1942] <= in[1138]; 
        out[1943] <= in[2588]; 
        out[1944] <= in[3567]; 
        out[1945] <= in[2510]; 
        out[1946] <= in[1634]; 
        out[1947] <= in[2378]; 
        out[1948] <= in[1080]; 
        out[1949] <= in[592]; 
        out[1950] <= in[611]; 
        out[1951] <= in[1318]; 
        out[1952] <= in[1053]; 
        out[1953] <= in[422]; 
        out[1954] <= in[702]; 
        out[1955] <= in[170]; 
        out[1956] <= in[1018]; 
        out[1957] <= in[727]; 
        out[1958] <= in[326]; 
        out[1959] <= in[2149]; 
        out[1960] <= in[1161]; 
        out[1961] <= in[638]; 
        out[1962] <= in[1193]; 
        out[1963] <= in[1790]; 
        out[1964] <= in[1066]; 
        out[1965] <= in[2576]; 
        out[1966] <= in[3667]; 
        out[1967] <= in[2176]; 
        out[1968] <= in[1092]; 
        out[1969] <= in[1948]; 
        out[1970] <= in[3806]; 
        out[1971] <= in[1441]; 
        out[1972] <= in[1788]; 
        out[1973] <= in[910]; 
        out[1974] <= in[2803]; 
        out[1975] <= in[1362]; 
        out[1976] <= in[820]; 
        out[1977] <= in[4094]; 
        out[1978] <= in[854]; 
        out[1979] <= in[46]; 
        out[1980] <= in[3543]; 
        out[1981] <= in[2263]; 
        out[1982] <= in[918]; 
        out[1983] <= in[3420]; 
        out[1984] <= in[3629]; 
        out[1985] <= in[413]; 
        out[1986] <= in[4057]; 
        out[1987] <= in[1040]; 
        out[1988] <= in[2391]; 
        out[1989] <= in[22]; 
        out[1990] <= in[3614]; 
        out[1991] <= in[1077]; 
        out[1992] <= in[2840]; 
        out[1993] <= in[3408]; 
        out[1994] <= in[2683]; 
        out[1995] <= in[3570]; 
        out[1996] <= in[3025]; 
        out[1997] <= in[2142]; 
        out[1998] <= in[429]; 
        out[1999] <= in[168]; 
        out[2000] <= in[196]; 
        out[2001] <= in[1323]; 
        out[2002] <= in[825]; 
        out[2003] <= in[3940]; 
        out[2004] <= in[515]; 
        out[2005] <= in[249]; 
        out[2006] <= in[319]; 
        out[2007] <= in[3073]; 
        out[2008] <= in[2711]; 
        out[2009] <= in[590]; 
        out[2010] <= in[3741]; 
        out[2011] <= in[38]; 
        out[2012] <= in[235]; 
        out[2013] <= in[1673]; 
        out[2014] <= in[3000]; 
        out[2015] <= in[3610]; 
        out[2016] <= in[3838]; 
        out[2017] <= in[2550]; 
        out[2018] <= in[3735]; 
        out[2019] <= in[3654]; 
        out[2020] <= in[2984]; 
        out[2021] <= in[478]; 
        out[2022] <= in[2442]; 
        out[2023] <= in[3613]; 
        out[2024] <= in[3747]; 
        out[2025] <= in[3799]; 
        out[2026] <= in[741]; 
        out[2027] <= in[4064]; 
        out[2028] <= in[2753]; 
        out[2029] <= in[1756]; 
        out[2030] <= in[469]; 
        out[2031] <= in[1864]; 
        out[2032] <= in[335]; 
        out[2033] <= in[1094]; 
        out[2034] <= in[3851]; 
        out[2035] <= in[2842]; 
        out[2036] <= in[3147]; 
        out[2037] <= in[839]; 
        out[2038] <= in[365]; 
        out[2039] <= in[4025]; 
        out[2040] <= in[4015]; 
        out[2041] <= in[3758]; 
        out[2042] <= in[954]; 
        out[2043] <= in[3832]; 
        out[2044] <= in[822]; 
        out[2045] <= in[3476]; 
        out[2046] <= in[1065]; 
        out[2047] <= in[1542]; 
        out[2048] <= in[3797]; 
        out[2049] <= in[1298]; 
        out[2050] <= in[311]; 
        out[2051] <= in[2204]; 
        out[2052] <= in[785]; 
        out[2053] <= in[1878]; 
        out[2054] <= in[118]; 
        out[2055] <= in[2272]; 
        out[2056] <= in[414]; 
        out[2057] <= in[2804]; 
        out[2058] <= in[1620]; 
        out[2059] <= in[3481]; 
        out[2060] <= in[2873]; 
        out[2061] <= in[2615]; 
        out[2062] <= in[1114]; 
        out[2063] <= in[3474]; 
        out[2064] <= in[1719]; 
        out[2065] <= in[3030]; 
        out[2066] <= in[3740]; 
        out[2067] <= in[3530]; 
        out[2068] <= in[2988]; 
        out[2069] <= in[1270]; 
        out[2070] <= in[817]; 
        out[2071] <= in[3944]; 
        out[2072] <= in[1916]; 
        out[2073] <= in[3710]; 
        out[2074] <= in[1852]; 
        out[2075] <= in[657]; 
        out[2076] <= in[72]; 
        out[2077] <= in[539]; 
        out[2078] <= in[2190]; 
        out[2079] <= in[1933]; 
        out[2080] <= in[3623]; 
        out[2081] <= in[4093]; 
        out[2082] <= in[1993]; 
        out[2083] <= in[136]; 
        out[2084] <= in[1036]; 
        out[2085] <= in[1446]; 
        out[2086] <= in[1969]; 
        out[2087] <= in[2858]; 
        out[2088] <= in[3714]; 
        out[2089] <= in[3997]; 
        out[2090] <= in[1285]; 
        out[2091] <= in[2630]; 
        out[2092] <= in[1912]; 
        out[2093] <= in[1811]; 
        out[2094] <= in[2813]; 
        out[2095] <= in[1135]; 
        out[2096] <= in[735]; 
        out[2097] <= in[3870]; 
        out[2098] <= in[1154]; 
        out[2099] <= in[661]; 
        out[2100] <= in[1029]; 
        out[2101] <= in[1845]; 
        out[2102] <= in[1017]; 
        out[2103] <= in[695]; 
        out[2104] <= in[1127]; 
        out[2105] <= in[3764]; 
        out[2106] <= in[1516]; 
        out[2107] <= in[2506]; 
        out[2108] <= in[790]; 
        out[2109] <= in[1850]; 
        out[2110] <= in[3829]; 
        out[2111] <= in[1434]; 
        out[2112] <= in[2910]; 
        out[2113] <= in[1428]; 
        out[2114] <= in[3591]; 
        out[2115] <= in[334]; 
        out[2116] <= in[3877]; 
        out[2117] <= in[3866]; 
        out[2118] <= in[3196]; 
        out[2119] <= in[540]; 
        out[2120] <= in[1491]; 
        out[2121] <= in[1866]; 
        out[2122] <= in[3071]; 
        out[2123] <= in[1333]; 
        out[2124] <= in[242]; 
        out[2125] <= in[1636]; 
        out[2126] <= in[884]; 
        out[2127] <= in[926]; 
        out[2128] <= in[1364]; 
        out[2129] <= in[1296]; 
        out[2130] <= in[271]; 
        out[2131] <= in[2181]; 
        out[2132] <= in[1520]; 
        out[2133] <= in[1465]; 
        out[2134] <= in[2423]; 
        out[2135] <= in[1245]; 
        out[2136] <= in[2195]; 
        out[2137] <= in[3998]; 
        out[2138] <= in[991]; 
        out[2139] <= in[3245]; 
        out[2140] <= in[3848]; 
        out[2141] <= in[942]; 
        out[2142] <= in[2341]; 
        out[2143] <= in[3676]; 
        out[2144] <= in[1813]; 
        out[2145] <= in[3528]; 
        out[2146] <= in[2780]; 
        out[2147] <= in[2949]; 
        out[2148] <= in[3631]; 
        out[2149] <= in[4074]; 
        out[2150] <= in[232]; 
        out[2151] <= in[2969]; 
        out[2152] <= in[2250]; 
        out[2153] <= in[3270]; 
        out[2154] <= in[1042]; 
        out[2155] <= in[3068]; 
        out[2156] <= in[3535]; 
        out[2157] <= in[2002]; 
        out[2158] <= in[2094]; 
        out[2159] <= in[3006]; 
        out[2160] <= in[646]; 
        out[2161] <= in[3136]; 
        out[2162] <= in[2718]; 
        out[2163] <= in[1531]; 
        out[2164] <= in[1390]; 
        out[2165] <= in[3142]; 
        out[2166] <= in[2688]; 
        out[2167] <= in[3106]; 
        out[2168] <= in[3276]; 
        out[2169] <= in[2426]; 
        out[2170] <= in[3324]; 
        out[2171] <= in[1433]; 
        out[2172] <= in[2412]; 
        out[2173] <= in[1849]; 
        out[2174] <= in[389]; 
        out[2175] <= in[3889]; 
        out[2176] <= in[668]; 
        out[2177] <= in[3634]; 
        out[2178] <= in[2465]; 
        out[2179] <= in[3887]; 
        out[2180] <= in[201]; 
        out[2181] <= in[1477]; 
        out[2182] <= in[301]; 
        out[2183] <= in[2668]; 
        out[2184] <= in[322]; 
        out[2185] <= in[3930]; 
        out[2186] <= in[3444]; 
        out[2187] <= in[222]; 
        out[2188] <= in[2849]; 
        out[2189] <= in[1601]; 
        out[2190] <= in[967]; 
        out[2191] <= in[3366]; 
        out[2192] <= in[550]; 
        out[2193] <= in[2372]; 
        out[2194] <= in[304]; 
        out[2195] <= in[775]; 
        out[2196] <= in[4021]; 
        out[2197] <= in[455]; 
        out[2198] <= in[2812]; 
        out[2199] <= in[4003]; 
        out[2200] <= in[1559]; 
        out[2201] <= in[2245]; 
        out[2202] <= in[2939]; 
        out[2203] <= in[2482]; 
        out[2204] <= in[913]; 
        out[2205] <= in[2243]; 
        out[2206] <= in[1049]; 
        out[2207] <= in[1100]; 
        out[2208] <= in[3669]; 
        out[2209] <= in[2597]; 
        out[2210] <= in[1211]; 
        out[2211] <= in[1985]; 
        out[2212] <= in[2763]; 
        out[2213] <= in[2119]; 
        out[2214] <= in[3316]; 
        out[2215] <= in[1139]; 
        out[2216] <= in[4066]; 
        out[2217] <= in[1988]; 
        out[2218] <= in[3519]; 
        out[2219] <= in[2179]; 
        out[2220] <= in[795]; 
        out[2221] <= in[2751]; 
        out[2222] <= in[961]; 
        out[2223] <= in[2327]; 
        out[2224] <= in[3096]; 
        out[2225] <= in[1807]; 
        out[2226] <= in[3742]; 
        out[2227] <= in[241]; 
        out[2228] <= in[488]; 
        out[2229] <= in[2862]; 
        out[2230] <= in[3088]; 
        out[2231] <= in[1194]; 
        out[2232] <= in[3988]; 
        out[2233] <= in[3215]; 
        out[2234] <= in[1151]; 
        out[2235] <= in[2875]; 
        out[2236] <= in[3240]; 
        out[2237] <= in[382]; 
        out[2238] <= in[3362]; 
        out[2239] <= in[3248]; 
        out[2240] <= in[793]; 
        out[2241] <= in[1936]; 
        out[2242] <= in[726]; 
        out[2243] <= in[633]; 
        out[2244] <= in[3730]; 
        out[2245] <= in[1947]; 
        out[2246] <= in[2725]; 
        out[2247] <= in[3494]; 
        out[2248] <= in[3057]; 
        out[2249] <= in[74]; 
        out[2250] <= in[561]; 
        out[2251] <= in[3678]; 
        out[2252] <= in[2505]; 
        out[2253] <= in[1931]; 
        out[2254] <= in[1885]; 
        out[2255] <= in[1271]; 
        out[2256] <= in[2031]; 
        out[2257] <= in[1558]; 
        out[2258] <= in[55]; 
        out[2259] <= in[3975]; 
        out[2260] <= in[2819]; 
        out[2261] <= in[364]; 
        out[2262] <= in[988]; 
        out[2263] <= in[3969]; 
        out[2264] <= in[351]; 
        out[2265] <= in[2595]; 
        out[2266] <= in[2186]; 
        out[2267] <= in[1297]; 
        out[2268] <= in[3754]; 
        out[2269] <= in[2866]; 
        out[2270] <= in[3849]; 
        out[2271] <= in[2951]; 
        out[2272] <= in[2107]; 
        out[2273] <= in[2408]; 
        out[2274] <= in[562]; 
        out[2275] <= in[2815]; 
        out[2276] <= in[903]; 
        out[2277] <= in[3228]; 
        out[2278] <= in[1530]; 
        out[2279] <= in[2769]; 
        out[2280] <= in[3636]; 
        out[2281] <= in[3067]; 
        out[2282] <= in[3341]; 
        out[2283] <= in[3271]; 
        out[2284] <= in[3588]; 
        out[2285] <= in[3112]; 
        out[2286] <= in[109]; 
        out[2287] <= in[341]; 
        out[2288] <= in[1301]; 
        out[2289] <= in[1728]; 
        out[2290] <= in[3552]; 
        out[2291] <= in[693]; 
        out[2292] <= in[1025]; 
        out[2293] <= in[3873]; 
        out[2294] <= in[3992]; 
        out[2295] <= in[3524]; 
        out[2296] <= in[754]; 
        out[2297] <= in[3012]; 
        out[2298] <= in[3618]; 
        out[2299] <= in[1732]; 
        out[2300] <= in[2621]; 
        out[2301] <= in[447]; 
        out[2302] <= in[3291]; 
        out[2303] <= in[2821]; 
        out[2304] <= in[1109]; 
        out[2305] <= in[740]; 
        out[2306] <= in[233]; 
        out[2307] <= in[2995]; 
        out[2308] <= in[3640]; 
        out[2309] <= in[767]; 
        out[2310] <= in[1048]; 
        out[2311] <= in[658]; 
        out[2312] <= in[3642]; 
        out[2313] <= in[2111]; 
        out[2314] <= in[4047]; 
        out[2315] <= in[730]; 
        out[2316] <= in[2212]; 
        out[2317] <= in[2788]; 
        out[2318] <= in[1625]; 
        out[2319] <= in[3344]; 
        out[2320] <= in[1287]; 
        out[2321] <= in[764]; 
        out[2322] <= in[970]; 
        out[2323] <= in[640]; 
        out[2324] <= in[3532]; 
        out[2325] <= in[1469]; 
        out[2326] <= in[464]; 
        out[2327] <= in[3231]; 
        out[2328] <= in[1699]; 
        out[2329] <= in[533]; 
        out[2330] <= in[1422]; 
        out[2331] <= in[3093]; 
        out[2332] <= in[1793]; 
        out[2333] <= in[3390]; 
        out[2334] <= in[1338]; 
        out[2335] <= in[670]; 
        out[2336] <= in[3061]; 
        out[2337] <= in[3554]; 
        out[2338] <= in[2568]; 
        out[2339] <= in[3568]; 
        out[2340] <= in[2253]; 
        out[2341] <= in[3156]; 
        out[2342] <= in[1197]; 
        out[2343] <= in[1817]; 
        out[2344] <= in[3630]; 
        out[2345] <= in[2635]; 
        out[2346] <= in[1904]; 
        out[2347] <= in[635]; 
        out[2348] <= in[2537]; 
        out[2349] <= in[315]; 
        out[2350] <= in[1233]; 
        out[2351] <= in[3198]; 
        out[2352] <= in[641]; 
        out[2353] <= in[2]; 
        out[2354] <= in[782]; 
        out[2355] <= in[188]; 
        out[2356] <= in[882]; 
        out[2357] <= in[2792]; 
        out[2358] <= in[3274]; 
        out[2359] <= in[1614]; 
        out[2360] <= in[3753]; 
        out[2361] <= in[483]; 
        out[2362] <= in[1322]; 
        out[2363] <= in[904]; 
        out[2364] <= in[3389]; 
        out[2365] <= in[3948]; 
        out[2366] <= in[9]; 
        out[2367] <= in[3157]; 
        out[2368] <= in[1789]; 
        out[2369] <= in[1294]; 
        out[2370] <= in[3478]; 
        out[2371] <= in[1707]; 
        out[2372] <= in[33]; 
        out[2373] <= in[1117]; 
        out[2374] <= in[1055]; 
        out[2375] <= in[1038]; 
        out[2376] <= in[1360]; 
        out[2377] <= in[2076]; 
        out[2378] <= in[76]; 
        out[2379] <= in[2219]; 
        out[2380] <= in[3105]; 
        out[2381] <= in[3616]; 
        out[2382] <= in[3840]; 
        out[2383] <= in[2404]; 
        out[2384] <= in[2102]; 
        out[2385] <= in[1714]; 
        out[2386] <= in[1940]; 
        out[2387] <= in[681]; 
        out[2388] <= in[3817]; 
        out[2389] <= in[2834]; 
        out[2390] <= in[2187]; 
        out[2391] <= in[3417]; 
        out[2392] <= in[1966]; 
        out[2393] <= in[617]; 
        out[2394] <= in[135]; 
        out[2395] <= in[2929]; 
        out[2396] <= in[3641]; 
        out[2397] <= in[739]; 
        out[2398] <= in[3350]; 
        out[2399] <= in[3117]; 
        out[2400] <= in[4026]; 
        out[2401] <= in[1896]; 
        out[2402] <= in[3283]; 
        out[2403] <= in[2990]; 
        out[2404] <= in[1412]; 
        out[2405] <= in[1923]; 
        out[2406] <= in[2337]; 
        out[2407] <= in[536]; 
        out[2408] <= in[2989]; 
        out[2409] <= in[501]; 
        out[2410] <= in[3382]; 
        out[2411] <= in[2610]; 
        out[2412] <= in[3748]; 
        out[2413] <= in[1598]; 
        out[2414] <= in[2126]; 
        out[2415] <= in[742]; 
        out[2416] <= in[2771]; 
        out[2417] <= in[325]; 
        out[2418] <= in[402]; 
        out[2419] <= in[2915]; 
        out[2420] <= in[3830]; 
        out[2421] <= in[688]; 
        out[2422] <= in[3562]; 
        out[2423] <= in[1561]; 
        out[2424] <= in[3752]; 
        out[2425] <= in[2940]; 
        out[2426] <= in[3759]; 
        out[2427] <= in[3193]; 
        out[2428] <= in[1421]; 
        out[2429] <= in[470]; 
        out[2430] <= in[3159]; 
        out[2431] <= in[2981]; 
        out[2432] <= in[2413]; 
        out[2433] <= in[95]; 
        out[2434] <= in[576]; 
        out[2435] <= in[250]; 
        out[2436] <= in[1072]; 
        out[2437] <= in[3426]; 
        out[2438] <= in[2775]; 
        out[2439] <= in[2169]; 
        out[2440] <= in[1840]; 
        out[2441] <= in[1599]; 
        out[2442] <= in[3454]; 
        out[2443] <= in[800]; 
        out[2444] <= in[2316]; 
        out[2445] <= in[2276]; 
        out[2446] <= in[733]; 
        out[2447] <= in[3512]; 
        out[2448] <= in[1043]; 
        out[2449] <= in[1951]; 
        out[2450] <= in[1078]; 
        out[2451] <= in[3751]; 
        out[2452] <= in[1669]; 
        out[2453] <= in[3804]; 
        out[2454] <= in[2140]; 
        out[2455] <= in[2491]; 
        out[2456] <= in[1889]; 
        out[2457] <= in[2654]; 
        out[2458] <= in[354]; 
        out[2459] <= in[474]; 
        out[2460] <= in[2520]; 
        out[2461] <= in[2396]; 
        out[2462] <= in[1405]; 
        out[2463] <= in[186]; 
        out[2464] <= in[2802]; 
        out[2465] <= in[3439]; 
        out[2466] <= in[1775]; 
        out[2467] <= in[2750]; 
        out[2468] <= in[1115]; 
        out[2469] <= in[91]; 
        out[2470] <= in[1189]; 
        out[2471] <= in[3110]; 
        out[2472] <= in[3151]; 
        out[2473] <= in[2628]; 
        out[2474] <= in[442]; 
        out[2475] <= in[221]; 
        out[2476] <= in[3277]; 
        out[2477] <= in[3691]; 
        out[2478] <= in[1637]; 
        out[2479] <= in[3937]; 
        out[2480] <= in[3312]; 
        out[2481] <= in[849]; 
        out[2482] <= in[1306]; 
        out[2483] <= in[2879]; 
        out[2484] <= in[566]; 
        out[2485] <= in[1274]; 
        out[2486] <= in[2447]; 
        out[2487] <= in[3845]; 
        out[2488] <= in[1820]; 
        out[2489] <= in[3138]; 
        out[2490] <= in[1663]; 
        out[2491] <= in[1064]; 
        out[2492] <= in[403]; 
        out[2493] <= in[1514]; 
        out[2494] <= in[2786]; 
        out[2495] <= in[4004]; 
        out[2496] <= in[445]; 
        out[2497] <= in[1455]; 
        out[2498] <= in[908]; 
        out[2499] <= in[34]; 
        out[2500] <= in[2474]; 
        out[2501] <= in[2618]; 
        out[2502] <= in[247]; 
        out[2503] <= in[2781]; 
        out[2504] <= in[282]; 
        out[2505] <= in[1501]; 
        out[2506] <= in[2598]; 
        out[2507] <= in[2039]; 
        out[2508] <= in[2808]; 
        out[2509] <= in[2220]; 
        out[2510] <= in[1074]; 
        out[2511] <= in[332]; 
        out[2512] <= in[814]; 
        out[2513] <= in[2869]; 
        out[2514] <= in[3860]; 
        out[2515] <= in[473]; 
        out[2516] <= in[3163]; 
        out[2517] <= in[2192]; 
        out[2518] <= in[680]; 
        out[2519] <= in[2052]; 
        out[2520] <= in[17]; 
        out[2521] <= in[1890]; 
        out[2522] <= in[1300]; 
        out[2523] <= in[3617]; 
        out[2524] <= in[3922]; 
        out[2525] <= in[768]; 
        out[2526] <= in[5]; 
        out[2527] <= in[165]; 
        out[2528] <= in[2943]; 
        out[2529] <= in[783]; 
        out[2530] <= in[2844]; 
        out[2531] <= in[2676]; 
        out[2532] <= in[794]; 
        out[2533] <= in[2852]; 
        out[2534] <= in[3503]; 
        out[2535] <= in[2138]; 
        out[2536] <= in[56]; 
        out[2537] <= in[284]; 
        out[2538] <= in[2226]; 
        out[2539] <= in[2757]; 
        out[2540] <= in[2544]; 
        out[2541] <= in[4065]; 
        out[2542] <= in[1972]; 
        out[2543] <= in[2726]; 
        out[2544] <= in[3226]; 
        out[2545] <= in[2100]; 
        out[2546] <= in[2766]; 
        out[2547] <= in[2870]; 
        out[2548] <= in[257]; 
        out[2549] <= in[456]; 
        out[2550] <= in[3831]; 
        out[2551] <= in[2000]; 
        out[2552] <= in[519]; 
        out[2553] <= in[2764]; 
        out[2554] <= in[2178]; 
        out[2555] <= in[2115]; 
        out[2556] <= in[2374]; 
        out[2557] <= in[3402]; 
        out[2558] <= in[3709]; 
        out[2559] <= in[3383]; 
        out[2560] <= in[3014]; 
        out[2561] <= in[1068]; 
        out[2562] <= in[2738]; 
        out[2563] <= in[3534]; 
        out[2564] <= in[3118]; 
        out[2565] <= in[3994]; 
        out[2566] <= in[1060]; 
        out[2567] <= in[2716]; 
        out[2568] <= in[1683]; 
        out[2569] <= in[3858]; 
        out[2570] <= in[923]; 
        out[2571] <= in[465]; 
        out[2572] <= in[3573]; 
        out[2573] <= in[2987]; 
        out[2574] <= in[1432]; 
        out[2575] <= in[683]; 
        out[2576] <= in[2483]; 
        out[2577] <= in[2469]; 
        out[2578] <= in[3202]; 
        out[2579] <= in[3569]; 
        out[2580] <= in[3416]; 
        out[2581] <= in[3078]; 
        out[2582] <= in[2589]; 
        out[2583] <= in[432]; 
        out[2584] <= in[1183]; 
        out[2585] <= in[1856]; 
        out[2586] <= in[2089]; 
        out[2587] <= in[3980]; 
        out[2588] <= in[1640]; 
        out[2589] <= in[430]; 
        out[2590] <= in[230]; 
        out[2591] <= in[3721]; 
        out[2592] <= in[3653]; 
        out[2593] <= in[718]; 
        out[2594] <= in[1213]; 
        out[2595] <= in[3210]; 
        out[2596] <= in[2651]; 
        out[2597] <= in[3098]; 
        out[2598] <= in[3409]; 
        out[2599] <= in[3486]; 
        out[2600] <= in[153]; 
        out[2601] <= in[24]; 
        out[2602] <= in[1005]; 
        out[2603] <= in[1198]; 
        out[2604] <= in[507]; 
        out[2605] <= in[3119]; 
        out[2606] <= in[3971]; 
        out[2607] <= in[3013]; 
        out[2608] <= in[394]; 
        out[2609] <= in[1009]; 
        out[2610] <= in[1687]; 
        out[2611] <= in[866]; 
        out[2612] <= in[2466]; 
        out[2613] <= in[3798]; 
        out[2614] <= in[180]; 
        out[2615] <= in[2136]; 
        out[2616] <= in[2425]; 
        out[2617] <= in[3619]; 
        out[2618] <= in[2768]; 
        out[2619] <= in[3356]; 
        out[2620] <= in[2043]; 
        out[2621] <= in[1968]; 
        out[2622] <= in[3328]; 
        out[2623] <= in[3820]; 
        out[2624] <= in[2567]; 
        out[2625] <= in[3578]; 
        out[2626] <= in[3368]; 
        out[2627] <= in[1861]; 
        out[2628] <= in[3459]; 
        out[2629] <= in[1453]; 
        out[2630] <= in[57]; 
        out[2631] <= in[1950]; 
        out[2632] <= in[1766]; 
        out[2633] <= in[1828]; 
        out[2634] <= in[2525]; 
        out[2635] <= in[3841]; 
        out[2636] <= in[4055]; 
        out[2637] <= in[757]; 
        out[2638] <= in[1868]; 
        out[2639] <= in[3325]; 
        out[2640] <= in[1886]; 
        out[2641] <= in[307]; 
        out[2642] <= in[573]; 
        out[2643] <= in[3546]; 
        out[2644] <= in[845]; 
        out[2645] <= in[669]; 
        out[2646] <= in[2746]; 
        out[2647] <= in[2496]; 
        out[2648] <= in[676]; 
        out[2649] <= in[1351]; 
        out[2650] <= in[2833]; 
        out[2651] <= in[2612]; 
        out[2652] <= in[431]; 
        out[2653] <= in[2501]; 
        out[2654] <= in[985]; 
        out[2655] <= in[1596]; 
        out[2656] <= in[2333]; 
        out[2657] <= in[2492]; 
        out[2658] <= in[3387]; 
        out[2659] <= in[1354]; 
        out[2660] <= in[3846]; 
        out[2661] <= in[3161]; 
        out[2662] <= in[3448]; 
        out[2663] <= in[821]; 
        out[2664] <= in[3954]; 
        out[2665] <= in[2246]; 
        out[2666] <= in[1510]; 
        out[2667] <= in[2933]; 
        out[2668] <= in[2968]; 
        out[2669] <= in[3066]; 
        out[2670] <= in[2397]; 
        out[2671] <= in[3192]; 
        out[2672] <= in[650]; 
        out[2673] <= in[1143]; 
        out[2674] <= in[2982]; 
        out[2675] <= in[2712]; 
        out[2676] <= in[579]; 
        out[2677] <= in[1622]; 
        out[2678] <= in[645]; 
        out[2679] <= in[2857]; 
        out[2680] <= in[243]; 
        out[2681] <= in[3001]; 
        out[2682] <= in[356]; 
        out[2683] <= in[3844]; 
        out[2684] <= in[3396]; 
        out[2685] <= in[45]; 
        out[2686] <= in[1436]; 
        out[2687] <= in[3525]; 
        out[2688] <= in[3559]; 
        out[2689] <= in[3265]; 
        out[2690] <= in[3209]; 
        out[2691] <= in[2605]; 
        out[2692] <= in[1946]; 
        out[2693] <= in[1123]; 
        out[2694] <= in[2168]; 
        out[2695] <= in[472]; 
        out[2696] <= in[2861]; 
        out[2697] <= in[1685]; 
        out[2698] <= in[691]; 
        out[2699] <= in[3133]; 
        out[2700] <= in[1922]; 
        out[2701] <= in[901]; 
        out[2702] <= in[1397]; 
        out[2703] <= in[3802]; 
        out[2704] <= in[434]; 
        out[2705] <= in[751]; 
        out[2706] <= in[2602]; 
        out[2707] <= in[517]; 
        out[2708] <= in[1677]; 
        out[2709] <= in[2158]; 
        out[2710] <= in[2349]; 
        out[2711] <= in[1202]; 
        out[2712] <= in[158]; 
        out[2713] <= in[1016]; 
        out[2714] <= in[2971]; 
        out[2715] <= in[1499]; 
        out[2716] <= in[832]; 
        out[2717] <= in[3626]; 
        out[2718] <= in[3990]; 
        out[2719] <= in[900]; 
        out[2720] <= in[925]; 
        out[2721] <= in[274]; 
        out[2722] <= in[1665]; 
        out[2723] <= in[555]; 
        out[2724] <= in[2649]; 
        out[2725] <= in[3908]; 
        out[2726] <= in[4020]; 
        out[2727] <= in[2009]; 
        out[2728] <= in[1130]; 
        out[2729] <= in[2432]; 
        out[2730] <= in[3290]; 
        out[2731] <= in[1050]; 
        out[2732] <= in[2614]; 
        out[2733] <= in[2922]; 
        out[2734] <= in[3144]; 
        out[2735] <= in[2173]; 
        out[2736] <= in[287]; 
        out[2737] <= in[117]; 
        out[2738] <= in[1552]; 
        out[2739] <= in[2153]; 
        out[2740] <= in[685]; 
        out[2741] <= in[2085]; 
        out[2742] <= in[762]; 
        out[2743] <= in[3520]; 
        out[2744] <= in[3373]; 
        out[2745] <= in[1462]; 
        out[2746] <= in[2268]; 
        out[2747] <= in[2511]; 
        out[2748] <= in[960]; 
        out[2749] <= in[3896]; 
        out[2750] <= in[1646]; 
        out[2751] <= in[88]; 
        out[2752] <= in[3991]; 
        out[2753] <= in[2291]; 
        out[2754] <= in[2065]; 
        out[2755] <= in[2859]; 
        out[2756] <= in[2662]; 
        out[2757] <= in[3973]; 
        out[2758] <= in[1125]; 
        out[2759] <= in[3483]; 
        out[2760] <= in[93]; 
        out[2761] <= in[1906]; 
        out[2762] <= in[605]; 
        out[2763] <= in[3650]; 
        out[2764] <= in[2381]; 
        out[2765] <= in[1429]; 
        out[2766] <= in[2051]; 
        out[2767] <= in[1502]; 
        out[2768] <= in[1228]; 
        out[2769] <= in[2837]; 
        out[2770] <= in[3601]; 
        out[2771] <= in[3043]; 
        out[2772] <= in[3207]; 
        out[2773] <= in[867]; 
        out[2774] <= in[2591]; 
        out[2775] <= in[3154]; 
        out[2776] <= in[1395]; 
        out[2777] <= in[328]; 
        out[2778] <= in[3060]; 
        out[2779] <= in[2344]; 
        out[2780] <= in[1774]; 
        out[2781] <= in[3645]; 
        out[2782] <= in[2827]; 
        out[2783] <= in[3146]; 
        out[2784] <= in[1391]; 
        out[2785] <= in[1486]; 
        out[2786] <= in[1546]; 
        out[2787] <= in[3440]; 
        out[2788] <= in[2818]; 
        out[2789] <= in[2562]; 
        out[2790] <= in[1444]; 
        out[2791] <= in[2486]; 
        out[2792] <= in[593]; 
        out[2793] <= in[3090]; 
        out[2794] <= in[883]; 
        out[2795] <= in[3256]; 
        out[2796] <= in[3475]; 
        out[2797] <= in[189]; 
        out[2798] <= in[1808]; 
        out[2799] <= in[132]; 
        out[2800] <= in[2955]; 
        out[2801] <= in[1862]; 
        out[2802] <= in[3783]; 
        out[2803] <= in[2384]; 
        out[2804] <= in[44]; 
        out[2805] <= in[752]; 
        out[2806] <= in[1515]; 
        out[2807] <= in[4071]; 
        out[2808] <= in[2906]; 
        out[2809] <= in[3865]; 
        out[2810] <= in[1905]; 
        out[2811] <= in[3477]; 
        out[2812] <= in[384]; 
        out[2813] <= in[1897]; 
        out[2814] <= in[1435]; 
        out[2815] <= in[859]; 
        out[2816] <= in[2160]; 
        out[2817] <= in[47]; 
        out[2818] <= in[4030]; 
        out[2819] <= in[1695]; 
        out[2820] <= in[3200]; 
        out[2821] <= in[672]; 
        out[2822] <= in[1483]; 
        out[2823] <= in[1141]; 
        out[2824] <= in[3549]; 
        out[2825] <= in[363]; 
        out[2826] <= in[4056]; 
        out[2827] <= in[387]; 
        out[2828] <= in[286]; 
        out[2829] <= in[2722]; 
        out[2830] <= in[3608]; 
        out[2831] <= in[41]; 
        out[2832] <= in[1738]; 
        out[2833] <= in[552]; 
        out[2834] <= in[1387]; 
        out[2835] <= in[3895]; 
        out[2836] <= in[2902]; 
        out[2837] <= in[83]; 
        out[2838] <= in[2117]; 
        out[2839] <= in[1260]; 
        out[2840] <= in[1780]; 
        out[2841] <= in[1859]; 
        out[2842] <= in[309]; 
        out[2843] <= in[613]; 
        out[2844] <= in[3508]; 
        out[2845] <= in[1099]; 
        out[2846] <= in[344]; 
        out[2847] <= in[870]; 
        out[2848] <= in[2817]; 
        out[2849] <= in[2001]; 
        out[2850] <= in[1875]; 
        out[2851] <= in[406]; 
        out[2852] <= in[1185]; 
        out[2853] <= in[2807]; 
        out[2854] <= in[2338]; 
        out[2855] <= in[804]; 
        out[2856] <= in[3695]; 
        out[2857] <= in[927]; 
        out[2858] <= in[1083]; 
        out[2859] <= in[1506]; 
        out[2860] <= in[2324]; 
        out[2861] <= in[1389]; 
        out[2862] <= in[3040]; 
        out[2863] <= in[268]; 
        out[2864] <= in[556]; 
        out[2865] <= in[1810]; 
        out[2866] <= in[1101]; 
        out[2867] <= in[824]; 
        out[2868] <= in[1666]; 
        out[2869] <= in[3258]; 
        out[2870] <= in[629]; 
        out[2871] <= in[2068]; 
        out[2872] <= in[1624]; 
        out[2873] <= in[2235]; 
        out[2874] <= in[2024]; 
        out[2875] <= in[2886]; 
        out[2876] <= in[3176]; 
        out[2877] <= in[3121]; 
        out[2878] <= in[3803]; 
        out[2879] <= in[2331]; 
        out[2880] <= in[3615]; 
        out[2881] <= in[29]; 
        out[2882] <= in[3072]; 
        out[2883] <= in[396]; 
        out[2884] <= in[2420]; 
        out[2885] <= in[529]; 
        out[2886] <= in[182]; 
        out[2887] <= in[4086]; 
        out[2888] <= in[3927]; 
        out[2889] <= in[1846]; 
        out[2890] <= in[2679]; 
        out[2891] <= in[3938]; 
        out[2892] <= in[3869]; 
        out[2893] <= in[276]; 
        out[2894] <= in[1703]; 
        out[2895] <= in[265]; 
        out[2896] <= in[921]; 
        out[2897] <= in[1407]; 
        out[2898] <= in[3850]; 
        out[2899] <= in[2180]; 
        out[2900] <= in[145]; 
        out[2901] <= in[1869]; 
        out[2902] <= in[3499]; 
        out[2903] <= in[1033]; 
        out[2904] <= in[2398]; 
        out[2905] <= in[1835]; 
        out[2906] <= in[3611]; 
        out[2907] <= in[375]; 
        out[2908] <= in[1388]; 
        out[2909] <= in[756]; 
        out[2910] <= in[3621]; 
        out[2911] <= in[3299]; 
        out[2912] <= in[997]; 
        out[2913] <= in[2062]; 
        out[2914] <= in[3398]; 
        out[2915] <= in[2957]; 
        out[2916] <= in[263]; 
        out[2917] <= in[2481]; 
        out[2918] <= in[841]; 
        out[2919] <= in[2619]; 
        out[2920] <= in[1063]; 
        out[2921] <= in[2144]; 
        out[2922] <= in[2351]; 
        out[2923] <= in[1524]; 
        out[2924] <= in[803]; 
        out[2925] <= in[549]; 
        out[2926] <= in[684]; 
        out[2927] <= in[202]; 
        out[2928] <= in[2003]; 
        out[2929] <= in[1733]; 
        out[2930] <= in[2228]; 
        out[2931] <= in[623]; 
        out[2932] <= in[1874]; 
        out[2933] <= in[2749]; 
        out[2934] <= in[706]; 
        out[2935] <= in[2278]; 
        out[2936] <= in[2185]; 
        out[2937] <= in[1639]; 
        out[2938] <= in[1574]; 
        out[2939] <= in[934]; 
        out[2940] <= in[2367]; 
        out[2941] <= in[320]; 
        out[2942] <= in[1070]; 
        out[2943] <= in[2429]; 
        out[2944] <= in[2044]; 
        out[2945] <= in[1313]; 
        out[2946] <= in[3005]; 
        out[2947] <= in[731]; 
        out[2948] <= in[2279]; 
        out[2949] <= in[66]; 
        out[2950] <= in[144]; 
        out[2951] <= in[1148]; 
        out[2952] <= in[2303]; 
        out[2953] <= in[2728]; 
        out[2954] <= in[844]; 
        out[2955] <= in[3315]; 
        out[2956] <= in[3750]; 
        out[2957] <= in[1302]; 
        out[2958] <= in[3900]; 
        out[2959] <= in[3232]; 
        out[2960] <= in[77]; 
        out[2961] <= in[802]; 
        out[2962] <= in[2717]; 
        out[2963] <= in[2304]; 
        out[2964] <= in[2867]; 
        out[2965] <= in[2267]; 
        out[2966] <= in[2574]; 
        out[2967] <= in[506]; 
        out[2968] <= in[1133]; 
        out[2969] <= in[3736]; 
        out[2970] <= in[3346]; 
        out[2971] <= in[272]; 
        out[2972] <= in[372]; 
        out[2973] <= in[788]; 
        out[2974] <= in[830]; 
        out[2975] <= in[1700]; 
        out[2976] <= in[3531]; 
        out[2977] <= in[2920]; 
        out[2978] <= in[2532]; 
        out[2979] <= in[3967]; 
        out[2980] <= in[1082]; 
        out[2981] <= in[1957]; 
        out[2982] <= in[1540]; 
        out[2983] <= in[3852]; 
        out[2984] <= in[2172]; 
        out[2985] <= in[496]; 
        out[2986] <= in[2067]; 
        out[2987] <= in[1335]; 
        out[2988] <= in[2247]; 
        out[2989] <= in[1680]; 
        out[2990] <= in[3612]; 
        out[2991] <= in[2199]; 
        out[2992] <= in[3719]; 
        out[2993] <= in[833]; 
        out[2994] <= in[468]; 
        out[2995] <= in[1246]; 
        out[2996] <= in[40]; 
        out[2997] <= in[1865]; 
        out[2998] <= in[2297]; 
        out[2999] <= in[3768]; 
        out[3000] <= in[2063]; 
        out[3001] <= in[608]; 
        out[3002] <= in[995]; 
        out[3003] <= in[1293]; 
        out[3004] <= in[2947]; 
        out[3005] <= in[2197]; 
        out[3006] <= in[2252]; 
        out[3007] <= in[15]; 
        out[3008] <= in[3330]; 
        out[3009] <= in[90]; 
        out[3010] <= in[2521]; 
        out[3011] <= in[1105]; 
        out[3012] <= in[120]; 
        out[3013] <= in[1734]; 
        out[3014] <= in[2463]; 
        out[3015] <= in[1276]; 
        out[3016] <= in[1226]; 
        out[3017] <= in[255]; 
        out[3018] <= in[3609]; 
        out[3019] <= in[171]; 
        out[3020] <= in[1560]; 
        out[3021] <= in[1482]; 
        out[3022] <= in[922]; 
        out[3023] <= in[2347]; 
        out[3024] <= in[3441]; 
        out[3025] <= in[39]; 
        out[3026] <= in[256]; 
        out[3027] <= in[678]; 
        out[3028] <= in[1674]; 
        out[3029] <= in[280]; 
        out[3030] <= in[2417]; 
        out[3031] <= in[197]; 
        out[3032] <= in[547]; 
        out[3033] <= in[3511]; 
        out[3034] <= in[330]; 
        out[3035] <= in[2691]; 
        out[3036] <= in[571]; 
        out[3037] <= in[2685]; 
        out[3038] <= in[4046]; 
        out[3039] <= in[1365]; 
        out[3040] <= in[3069]; 
        out[3041] <= in[1363]; 
        out[3042] <= in[3996]; 
        out[3043] <= in[2129]; 
        out[3044] <= in[3594]; 
        out[3045] <= in[1314]; 
        out[3046] <= in[2918]; 
        out[3047] <= in[4019]; 
        out[3048] <= in[1106]; 
        out[3049] <= in[3137]; 
        out[3050] <= in[191]; 
        out[3051] <= in[1980]; 
        out[3052] <= in[3051]; 
        out[3053] <= in[2493]; 
        out[3054] <= in[3303]; 
        out[3055] <= in[2664]; 
        out[3056] <= in[1583]; 
        out[3057] <= in[842]; 
        out[3058] <= in[2106]; 
        out[3059] <= in[2459]; 
        out[3060] <= in[2911]; 
        out[3061] <= in[2904]; 
        out[3062] <= in[267]; 
        out[3063] <= in[3230]; 
        out[3064] <= in[2958]; 
        out[3065] <= in[1403]; 
        out[3066] <= in[1585]; 
        out[3067] <= in[3956]; 
        out[3068] <= in[3715]; 
        out[3069] <= in[2609]; 
        out[3070] <= in[1976]; 
        out[3071] <= in[624]; 
        out[3072] <= in[3491]; 
        out[3073] <= in[2071]; 
        out[3074] <= in[3213]; 
        out[3075] <= in[374]; 
        out[3076] <= in[3705]; 
        out[3077] <= in[935]; 
        out[3078] <= in[2021]; 
        out[3079] <= in[3504]; 
        out[3080] <= in[919]; 
        out[3081] <= in[2450]; 
        out[3082] <= in[2213]; 
        out[3083] <= in[3769]; 
        out[3084] <= in[3995]; 
        out[3085] <= in[2323]; 
        out[3086] <= in[3445]; 
        out[3087] <= in[2175]; 
        out[3088] <= in[1352]; 
        out[3089] <= in[1653]; 
        out[3090] <= in[1445]; 
        out[3091] <= in[697]; 
        out[3092] <= in[909]; 
        out[3093] <= in[992]; 
        out[3094] <= in[2707]; 
        out[3095] <= in[916]; 
        out[3096] <= in[42]; 
        out[3097] <= in[3313]; 
        out[3098] <= in[2992]; 
        out[3099] <= in[732]; 
        out[3100] <= in[3909]; 
        out[3101] <= in[1611]; 
        out[3102] <= in[3250]; 
        out[3103] <= in[1305]; 
        out[3104] <= in[2850]; 
        out[3105] <= in[1203]; 
        out[3106] <= in[2154]; 
        out[3107] <= in[1851]; 
        out[3108] <= in[2694]; 
        out[3109] <= in[1309]; 
        out[3110] <= in[2234]; 
        out[3111] <= in[1508]; 
        out[3112] <= in[2358]; 
        out[3113] <= in[2549]; 
        out[3114] <= in[3095]; 
        out[3115] <= in[1782]; 
        out[3116] <= in[420]; 
        out[3117] <= in[3514]; 
        out[3118] <= in[1373]; 
        out[3119] <= in[2556]; 
        out[3120] <= in[1111]; 
        out[3121] <= in[415]; 
        out[3122] <= in[1659]; 
        out[3123] <= in[952]; 
        out[3124] <= in[920]; 
        out[3125] <= in[3431]; 
        out[3126] <= in[3718]; 
        out[3127] <= in[3796]; 
        out[3128] <= in[2644]; 
        out[3129] <= in[2269]; 
        out[3130] <= in[580]; 
        out[3131] <= in[1085]; 
        out[3132] <= in[3285]; 
        out[3133] <= in[291]; 
        out[3134] <= in[398]; 
        out[3135] <= in[2845]; 
        out[3136] <= in[1348]; 
        out[3137] <= in[3334]; 
        out[3138] <= in[587]; 
        out[3139] <= in[545]; 
        out[3140] <= in[1761]; 
        out[3141] <= in[3395]; 
        out[3142] <= in[2891]; 
        out[3143] <= in[3711]; 
        out[3144] <= in[3089]; 
        out[3145] <= in[664]; 
        out[3146] <= in[1084]; 
        out[3147] <= in[696]; 
        out[3148] <= in[1142]; 
        out[3149] <= in[1457]; 
        out[3150] <= in[175]; 
        out[3151] <= in[361]; 
        out[3152] <= in[3731]; 
        out[3153] <= in[3679]; 
        out[3154] <= in[987]; 
        out[3155] <= in[1967]; 
        out[3156] <= in[3538]; 
        out[3157] <= in[3970]; 
        out[3158] <= in[1047]; 
        out[3159] <= in[3781]; 
        out[3160] <= in[1345]; 
        out[3161] <= in[3732]; 
        out[3162] <= in[503]; 
        out[3163] <= in[3049]; 
        out[3164] <= in[96]; 
        out[3165] <= in[2742]; 
        out[3166] <= in[3502]; 
        out[3167] <= in[4034]; 
        out[3168] <= in[3770]; 
        out[3169] <= in[1855]; 
        out[3170] <= in[3460]; 
        out[3171] <= in[1652]; 
        out[3172] <= in[1900]; 
        out[3173] <= in[1643]; 
        out[3174] <= in[3648]; 
        out[3175] <= in[300]; 
        out[3176] <= in[3086]; 
        out[3177] <= in[3041]; 
        out[3178] <= in[4001]; 
        out[3179] <= in[801]; 
        out[3180] <= in[2830]; 
        out[3181] <= in[781]; 
        out[3182] <= in[1031]; 
        out[3183] <= in[3430]; 
        out[3184] <= in[4039]; 
        out[3185] <= in[4038]; 
        out[3186] <= in[3652]; 
        out[3187] <= in[1716]; 
        out[3188] <= in[2572]; 
        out[3189] <= in[1447]; 
        out[3190] <= in[779]; 
        out[3191] <= in[3668]; 
        out[3192] <= in[2795]; 
        out[3193] <= in[3488]; 
        out[3194] <= in[495]; 
        out[3195] <= in[1396]; 
        out[3196] <= in[3288]; 
        out[3197] <= in[686]; 
        out[3198] <= in[1088]; 
        out[3199] <= in[3314]; 
        out[3200] <= in[2435]; 
        out[3201] <= in[933]; 
        out[3202] <= in[369]; 
        out[3203] <= in[1410]; 
        out[3204] <= in[3279]; 
        out[3205] <= in[1369]; 
        out[3206] <= in[1672]; 
        out[3207] <= in[3907]; 
        out[3208] <= in[218]; 
        out[3209] <= in[2670]; 
        out[3210] <= in[1116]; 
        out[3211] <= in[3697]; 
        out[3212] <= in[3893]; 
        out[3213] <= in[1978]; 
        out[3214] <= in[3941]; 
        out[3215] <= in[1140]; 
        out[3216] <= in[504]; 
        out[3217] <= in[43]; 
        out[3218] <= in[318]; 
        out[3219] <= in[936]; 
        out[3220] <= in[89]; 
        out[3221] <= in[80]; 
        out[3222] <= in[1954]; 
        out[3223] <= in[1908]; 
        out[3224] <= in[3681]; 
        out[3225] <= in[891]; 
        out[3226] <= in[710]; 
        out[3227] <= in[70]; 
        out[3228] <= in[2974]; 
        out[3229] <= in[1252]; 
        out[3230] <= in[707]; 
        out[3231] <= in[3763]; 
        out[3232] <= in[3487]; 
        out[3233] <= in[4000]; 
        out[3234] <= in[1171]; 
        out[3235] <= in[324]; 
        out[3236] <= in[3463]; 
        out[3237] <= in[2345]; 
        out[3238] <= in[1602]; 
        out[3239] <= in[2336]; 
        out[3240] <= in[947]; 
        out[3241] <= in[1592]; 
        out[3242] <= in[979]; 
        out[3243] <= in[1576]; 
        out[3244] <= in[2893]; 
        out[3245] <= in[1577]; 
        out[3246] <= in[2132]; 
        out[3247] <= in[1230]; 
        out[3248] <= in[3167]; 
        out[3249] <= in[912]; 
        out[3250] <= in[1983]; 
        out[3251] <= in[3436]; 
        out[3252] <= in[1058]; 
        out[3253] <= in[1500]; 
        out[3254] <= in[3815]; 
        out[3255] <= in[760]; 
        out[3256] <= in[106]; 
        out[3257] <= in[2048]; 
        out[3258] <= in[2701]; 
        out[3259] <= in[3649]; 
        out[3260] <= in[2629]; 
        out[3261] <= in[1741]; 
        out[3262] <= in[2710]; 
        out[3263] <= in[690]; 
        out[3264] <= in[62]; 
        out[3265] <= in[1474]; 
        out[3266] <= in[853]; 
        out[3267] <= in[2695]; 
        out[3268] <= in[1537]; 
        out[3269] <= in[2242]; 
        out[3270] <= in[19]; 
        out[3271] <= in[3664]; 
        out[3272] <= in[2998]; 
        out[3273] <= in[1218]; 
        out[3274] <= in[2983]; 
        out[3275] <= in[240]; 
        out[3276] <= in[1754]; 
        out[3277] <= in[67]; 
        out[3278] <= in[2237]; 
        out[3279] <= in[3393]; 
        out[3280] <= in[1584]; 
        out[3281] <= in[772]; 
        out[3282] <= in[1839]; 
        out[3283] <= in[1201]; 
        out[3284] <= in[3836]; 
        out[3285] <= in[2953]; 
        out[3286] <= in[4024]; 
        out[3287] <= in[2034]; 
        out[3288] <= in[2162]; 
        out[3289] <= in[1854]; 
        out[3290] <= in[3323]; 
        out[3291] <= in[1071]; 
        out[3292] <= in[2785]; 
        out[3293] <= in[2339]; 
        out[3294] <= in[1006]; 
        out[3295] <= in[1694]; 
        out[3296] <= in[1272]; 
        out[3297] <= in[2674]; 
        out[3298] <= in[449]; 
        out[3299] <= in[125]; 
        out[3300] <= in[1538]; 
        out[3301] <= in[423]; 
        out[3302] <= in[3241]; 
        out[3303] <= in[546]; 
        out[3304] <= in[994]; 
        out[3305] <= in[2836]; 
        out[3306] <= in[3199]; 
        out[3307] <= in[1236]; 
        out[3308] <= in[1724]; 
        out[3309] <= in[2607]; 
        out[3310] <= in[2112]; 
        out[3311] <= in[616]; 
        out[3312] <= in[1167]; 
        out[3313] <= in[1209]; 
        out[3314] <= in[3470]; 
        out[3315] <= in[747]; 
        out[3316] <= in[930]; 
        out[3317] <= in[2648]; 
        out[3318] <= in[2191]; 
        out[3319] <= in[1629]; 
        out[3320] <= in[1648]; 
        out[3321] <= in[283]; 
        out[3322] <= in[3217]; 
        out[3323] <= in[2040]; 
        out[3324] <= in[3472]; 
        out[3325] <= in[486]; 
        out[3326] <= in[1956]; 
        out[3327] <= in[3565]; 
        out[3328] <= in[876]; 
        out[3329] <= in[2671]; 
        out[3330] <= in[3065]; 
        out[3331] <= in[2332]; 
        out[3332] <= in[2352]; 
        out[3333] <= in[1942]; 
        out[3334] <= in[911]; 
        out[3335] <= in[1013]; 
        out[3336] <= in[1319]; 
        out[3337] <= in[81]; 
        out[3338] <= in[755]; 
        out[3339] <= in[298]; 
        out[3340] <= in[1876]; 
        out[3341] <= in[3224]; 
        out[3342] <= in[1631]; 
        out[3343] <= in[2673]; 
        out[3344] <= in[3165]; 
        out[3345] <= in[1910]; 
        out[3346] <= in[4029]; 
        out[3347] <= in[1926]; 
        out[3348] <= in[3269]; 
        out[3349] <= in[2762]; 
        out[3350] <= in[3910]; 
        out[3351] <= in[3195]; 
        out[3352] <= in[1713]; 
        out[3353] <= in[2560]; 
        out[3354] <= in[3964]; 
        out[3355] <= in[701]; 
        out[3356] <= in[3406]; 
        out[3357] <= in[225]; 
        out[3358] <= in[3259]; 
        out[3359] <= in[3729]; 
        out[3360] <= in[1752]; 
        out[3361] <= in[21]; 
        out[3362] <= in[2334]; 
        out[3363] <= in[2320]; 
        out[3364] <= in[3082]; 
        out[3365] <= in[2706]; 
        out[3366] <= in[1964]; 
        out[3367] <= in[522]; 
        out[3368] <= in[3946]; 
        out[3369] <= in[3188]; 
        out[3370] <= in[774]; 
        out[3371] <= in[850]; 
        out[3372] <= in[3120]; 
        out[3373] <= in[494]; 
        out[3374] <= in[1149]; 
        out[3375] <= in[2399]; 
        out[3376] <= in[3550]; 
        out[3377] <= in[302]; 
        out[3378] <= in[3928]; 
        out[3379] <= in[1254]; 
        out[3380] <= in[2714]; 
        out[3381] <= in[2177]; 
        out[3382] <= in[1113]; 
        out[3383] <= in[2066]; 
        out[3384] <= in[3085]; 
        out[3385] <= in[597]; 
        out[3386] <= in[1350]; 
        out[3387] <= in[1431]; 
        out[3388] <= in[1174]; 
        out[3389] <= in[1458]; 
        out[3390] <= in[2203]; 
        out[3391] <= in[1860]; 
        out[3392] <= in[1986]; 
        out[3393] <= in[2594]; 
        out[3394] <= in[20]; 
        out[3395] <= in[2512]; 
        out[3396] <= in[137]; 
        out[3397] <= in[279]; 
        out[3398] <= in[1818]; 
        out[3399] <= in[964]; 
        out[3400] <= in[600]; 
        out[3401] <= in[2854]; 
        out[3402] <= in[3987]; 
        out[3403] <= in[3541]; 
        out[3404] <= in[3026]; 
        out[3405] <= in[373]; 
        out[3406] <= in[940]; 
        out[3407] <= in[2699]; 
        out[3408] <= in[1579]; 
        out[3409] <= in[1824]; 
        out[3410] <= in[2361]; 
        out[3411] <= in[1164]; 
        out[3412] <= in[1108]; 
        out[3413] <= in[1359]; 
        out[3414] <= in[1772]; 
        out[3415] <= in[1487]; 
        out[3416] <= in[2265]; 
        out[3417] <= in[3521]; 
        out[3418] <= in[2523]; 
        out[3419] <= in[2084]; 
        out[3420] <= in[2141]; 
        out[3421] <= in[2799]; 
        out[3422] <= in[4075]; 
        out[3423] <= in[65]; 
        out[3424] <= in[116]; 
        out[3425] <= in[3963]; 
        out[3426] <= in[3694]; 
        out[3427] <= in[3911]; 
        out[3428] <= in[2801]; 
        out[3429] <= in[1831]; 
        out[3430] <= in[2543]; 
        out[3431] <= in[1004]; 
        out[3432] <= in[3469]; 
        out[3433] <= in[1909]; 
        out[3434] <= in[2161]; 
        out[3435] <= in[3242]; 
        out[3436] <= in[1797]; 
        out[3437] <= in[1181]; 
        out[3438] <= in[1726]; 
        out[3439] <= in[3789]; 
        out[3440] <= in[1103]; 
        out[3441] <= in[548]; 
        out[3442] <= in[2774]; 
        out[3443] <= in[3542]; 
        out[3444] <= in[2914]; 
        out[3445] <= in[3899]; 
        out[3446] <= in[1873]; 
        out[3447] <= in[3351]; 
        out[3448] <= in[1901]; 
        out[3449] <= in[3767]; 
        out[3450] <= in[719]; 
        out[3451] <= in[2330]; 
        out[3452] <= in[194]; 
        out[3453] <= in[888]; 
        out[3454] <= in[560]; 
        out[3455] <= in[750]; 
        out[3456] <= in[3304]; 
        out[3457] <= in[2468]; 
        out[3458] <= in[3391]; 
        out[3459] <= in[3771]; 
        out[3460] <= in[1091]; 
        out[3461] <= in[2462]; 
        out[3462] <= in[823]; 
        out[3463] <= in[3746]; 
        out[3464] <= in[3164]; 
        out[3465] <= in[2905]; 
        out[3466] <= in[3160]; 
        out[3467] <= in[984]; 
        out[3468] <= in[3662]; 
        out[3469] <= in[1792]; 
        out[3470] <= in[1470]; 
        out[3471] <= in[3319]; 
        out[3472] <= in[333]; 
        out[3473] <= in[3677]; 
        out[3474] <= in[2231]; 
        out[3475] <= in[1081]; 
        out[3476] <= in[1548]; 
        out[3477] <= in[2945]; 
        out[3478] <= in[448]; 
        out[3479] <= in[2007]; 
        out[3480] <= in[1182]; 
        out[3481] <= in[1773]; 
        out[3482] <= in[1291]; 
        out[3483] <= in[1485]; 
        out[3484] <= in[2047]; 
        out[3485] <= in[1880]; 
        out[3486] <= in[2497]; 
        out[3487] <= in[1881]; 
        out[3488] <= in[3297]; 
        out[3489] <= in[1693]; 
        out[3490] <= in[3361]; 
        out[3491] <= in[3882]; 
        out[3492] <= in[371]; 
        out[3493] <= in[1366]; 
        out[3494] <= in[542]; 
        out[3495] <= in[3172]; 
        out[3496] <= in[766]; 
        out[3497] <= in[3360]; 
        out[3498] <= in[1664]; 
        out[3499] <= in[3923]; 
        out[3500] <= in[3881]; 
        out[3501] <= in[1095]; 
        out[3502] <= in[1324]; 
        out[3503] <= in[1594]; 
        out[3504] <= in[2386]; 
        out[3505] <= in[738]; 
        out[3506] <= in[103]; 
        out[3507] <= in[3397]; 
        out[3508] <= in[3863]; 
        out[3509] <= in[2101]; 
        out[3510] <= in[3171]; 
        out[3511] <= in[337]; 
        out[3512] <= in[3926]; 
        out[3513] <= in[71]; 
        out[3514] <= in[79]; 
        out[3515] <= in[1155]; 
        out[3516] <= in[3600]; 
        out[3517] <= in[451]; 
        out[3518] <= in[208]; 
        out[3519] <= in[3773]; 
        out[3520] <= in[846]; 
        out[3521] <= in[873]; 
        out[3522] <= in[3665]; 
        out[3523] <= in[3760]; 
        out[3524] <= in[2569]; 
        out[3525] <= in[407]; 
        out[3526] <= in[2287]; 
        out[3527] <= in[1635]; 
        out[3528] <= in[2127]; 
        out[3529] <= in[1955]; 
        out[3530] <= in[1205]; 
        out[3531] <= in[1035]; 
        out[3532] <= in[1427]; 
        out[3533] <= in[989]; 
        out[3534] <= in[142]; 
        out[3535] <= in[2600]; 
        out[3536] <= in[462]; 
        out[3537] <= in[3620]; 
        out[3538] <= in[1841]; 
        out[3539] <= in[1124]; 
        out[3540] <= in[2033]; 
        out[3541] <= in[2965]; 
        out[3542] <= in[2022]; 
        out[3543] <= in[348]; 
        out[3544] <= in[485]; 
        out[3545] <= in[3933]; 
        out[3546] <= in[2097]; 
        out[3547] <= in[454]; 
        out[3548] <= in[18]; 
        out[3549] <= in[2035]; 
        out[3550] <= in[2359]; 
        out[3551] <= in[1762]; 
        out[3552] <= in[1120]; 
        out[3553] <= in[110]; 
        out[3554] <= in[1932]; 
        out[3555] <= in[2294]; 
        out[3556] <= in[1984]; 
        out[3557] <= in[843]; 
        out[3558] <= in[3777]; 
        out[3559] <= in[810]; 
        out[3560] <= in[1770]; 
        out[3561] <= in[559]; 
        out[3562] <= in[692]; 
        out[3563] <= in[2727]; 
        out[3564] <= in[147]; 
        out[3565] <= in[1089]; 
        out[3566] <= in[744]; 
        out[3567] <= in[3936]; 
        out[3568] <= in[49]; 
        out[3569] <= in[404]; 
        out[3570] <= in[316]; 
        out[3571] <= in[610]; 
        out[3572] <= in[558]; 
        out[3573] <= in[2991]; 
        out[3574] <= in[1580]; 
        out[3575] <= in[4040]; 
        out[3576] <= in[98]; 
        out[3577] <= in[2729]; 
        out[3578] <= in[1449]; 
        out[3579] <= in[2620]; 
        out[3580] <= in[2631]; 
        out[3581] <= in[1795]; 
        out[3582] <= in[2778]; 
        out[3583] <= in[713]; 
        out[3584] <= in[4006]; 
        out[3585] <= in[1172]; 
        out[3586] <= in[1002]; 
        out[3587] <= in[2900]; 
        out[3588] <= in[2049]; 
        out[3589] <= in[2564]; 
        out[3590] <= in[3329]; 
        out[3591] <= in[813]; 
        out[3592] <= in[126]; 
        out[3593] <= in[2064]; 
        out[3594] <= in[1837]; 
        out[3595] <= in[2700]; 
        out[3596] <= in[2926]; 
        out[3597] <= in[2414]; 
        out[3598] <= in[2793]; 
        out[3599] <= in[578]; 
        out[3600] <= in[2724]; 
        out[3601] <= in[1991]; 
        out[3602] <= in[2584]; 
        out[3603] <= in[1384]; 
        out[3604] <= in[3972]; 
        out[3605] <= in[3442]; 
        out[3606] <= in[4054]; 
        out[3607] <= in[2251]; 
        out[3608] <= in[3589]; 
        out[3609] <= in[308]; 
        out[3610] <= in[1096]; 
        out[3611] <= in[1533]; 
        out[3612] <= in[2312]; 
        out[3613] <= in[2053]; 
        out[3614] <= in[567]; 
        out[3615] <= in[784]; 
        out[3616] <= in[3177]; 
        out[3617] <= in[2585]; 
        out[3618] <= in[2883]; 
        out[3619] <= in[2166]; 
        out[3620] <= in[3145]; 
        out[3621] <= in[3485]; 
        out[3622] <= in[570]; 
        out[3623] <= in[2322]; 
        out[3624] <= in[1337]; 
        out[3625] <= in[3298]; 
        out[3626] <= in[4089]; 
        out[3627] <= in[2433]; 
        out[3628] <= in[3462]; 
        out[3629] <= in[498]; 
        out[3630] <= in[2494]; 
        out[3631] <= in[2765]; 
        out[3632] <= in[4088]; 
        out[3633] <= in[3002]; 
        out[3634] <= in[2865]; 
        out[3635] <= in[1383]; 
        out[3636] <= in[2418]; 
        out[3637] <= in[2657]; 
        out[3638] <= in[2202]; 
        out[3639] <= in[2503]; 
        out[3640] <= in[652]; 
        out[3641] <= in[3606]; 
        out[3642] <= in[1032]; 
        out[3643] <= in[1745]; 
        out[3644] <= in[346]; 
        out[3645] <= in[2449]; 
        out[3646] <= in[3204]; 
        out[3647] <= in[452]; 
        out[3648] <= in[724]; 
        out[3649] <= in[2596]; 
        out[3650] <= in[3301]; 
        out[3651] <= in[1982]; 
        out[3652] <= in[2528]; 
        out[3653] <= in[3257]; 
        out[3654] <= in[3599]; 
        out[3655] <= in[2309]; 
        out[3656] <= in[105]; 
        out[3657] <= in[3428]; 
        out[3658] <= in[2913]; 
        out[3659] <= in[59]; 
        out[3660] <= in[3810]; 
        out[3661] <= in[3208]; 
        out[3662] <= in[2809]; 
        out[3663] <= in[2709]; 
        out[3664] <= in[1424]; 
        out[3665] <= in[2114]; 
        out[3666] <= in[568]; 
        out[3667] <= in[3510]; 
        out[3668] <= in[78]; 
        out[3669] <= in[2055]; 
        out[3670] <= in[3019]; 
        out[3671] <= in[2379]; 
        out[3672] <= in[932]; 
        out[3673] <= in[2411]; 
        out[3674] <= in[2441]; 
        out[3675] <= in[2708]; 
        out[3676] <= in[1372]; 
        out[3677] <= in[383]; 
        out[3678] <= in[2603]; 
        out[3679] <= in[4033]; 
        out[3680] <= in[3353]; 
        out[3681] <= in[2782]; 
        out[3682] <= in[385]; 
        out[3683] <= in[3507]; 
        out[3684] <= in[2623]; 
        out[3685] <= in[3955]; 
        out[3686] <= in[3670]; 
        out[3687] <= in[639]; 
        out[3688] <= in[2125]; 
        out[3689] <= in[26]; 
        out[3690] <= in[2428]; 
        out[3691] <= in[2293]; 
        out[3692] <= in[3774]; 
        out[3693] <= in[3126]; 
        out[3694] <= in[1783]; 
        out[3695] <= in[3657]; 
        out[3696] <= in[3914]; 
        out[3697] <= in[3045]; 
        out[3698] <= in[1340]; 
        out[3699] <= in[60]; 
        out[3700] <= in[2977]; 
        out[3701] <= in[1570]; 
        out[3702] <= in[3780]; 
        out[3703] <= in[3989]; 
        out[3704] <= in[2453]; 
        out[3705] <= in[2407]; 
        out[3706] <= in[1825]; 
        out[3707] <= in[1504]; 
        out[3708] <= in[1877]; 
        out[3709] <= in[127]; 
        out[3710] <= in[1180]; 
        out[3711] <= in[1234]; 
        out[3712] <= in[3348]; 
        out[3713] <= in[1227]; 
        out[3714] <= in[872]; 
        out[3715] <= in[262]; 
        out[3716] <= in[2864]; 
        out[3717] <= in[2155]; 
        out[3718] <= in[3738]; 
        out[3719] <= in[2529]; 
        out[3720] <= in[295]; 
        out[3721] <= in[2388]; 
        out[3722] <= in[489]; 
        out[3723] <= in[2748]; 
        out[3724] <= in[2394]; 
        out[3725] <= in[1037]; 
        out[3726] <= in[1200]; 
        out[3727] <= in[1822]; 
        out[3728] <= in[435]; 
        out[3729] <= in[163]; 
        out[3730] <= in[1578]; 
        out[3731] <= in[416]; 
        out[3732] <= in[3223]; 
        out[3733] <= in[1057]; 
        out[3734] <= in[787]; 
        out[3735] <= in[2020]; 
        out[3736] <= in[2210]; 
        out[3737] <= in[3174]; 
        out[3738] <= in[728]; 
        out[3739] <= in[1232]; 
        out[3740] <= in[3044]; 
        out[3741] <= in[3544]; 
        out[3742] <= in[2262]; 
        out[3743] <= in[2740]; 
        out[3744] <= in[377]; 
        out[3745] <= in[1217]; 
        out[3746] <= in[881]; 
        out[3747] <= in[1943]; 
        out[3748] <= in[1269]; 
        out[3749] <= in[1019]; 
        out[3750] <= in[4061]; 
        out[3751] <= in[2997]; 
        out[3752] <= in[1573]; 
        out[3753] <= in[950]; 
        out[3754] <= in[835]; 
        out[3755] <= in[3813]; 
        out[3756] <= in[1834]; 
        out[3757] <= in[3132]; 
        out[3758] <= in[209]; 
        out[3759] <= in[1785]; 
        out[3760] <= in[1844]; 
        out[3761] <= in[655]; 
        out[3762] <= in[2994]; 
        out[3763] <= in[1231]; 
        out[3764] <= in[1408]; 
        out[3765] <= in[2029]; 
        out[3766] <= in[3064]; 
        out[3767] <= in[4069]; 
        out[3768] <= in[1507]; 
        out[3769] <= in[2189]; 
        out[3770] <= in[3915]; 
        out[3771] <= in[2601]; 
        out[3772] <= in[2124]; 
        out[3773] <= in[261]; 
        out[3774] <= in[3447]; 
        out[3775] <= in[4090]; 
        out[3776] <= in[860]; 
        out[3777] <= in[2954]; 
        out[3778] <= in[2288]; 
        out[3779] <= in[2393]; 
        out[3780] <= in[1443]; 
        out[3781] <= in[1400]; 
        out[3782] <= in[1196]; 
        out[3783] <= in[1705]; 
        out[3784] <= in[1104]; 
        out[3785] <= in[2123]; 
        out[3786] <= in[3833]; 
        out[3787] <= in[945]; 
        out[3788] <= in[3206]; 
        out[3789] <= in[1809]; 
        out[3790] <= in[4077]; 
        out[3791] <= in[1425]; 
        out[3792] <= in[3131]; 
        out[3793] <= in[3560]; 
        out[3794] <= in[2580]; 
        out[3795] <= in[3722]; 
        out[3796] <= in[359]; 
        out[3797] <= in[3233]; 
        out[3798] <= in[2238]; 
        out[3799] <= in[2626]; 
        out[3800] <= in[2354]; 
        out[3801] <= in[553]; 
        out[3802] <= in[289]; 
        out[3803] <= in[588]; 
        out[3804] <= in[329]; 
        out[3805] <= in[1152]; 
        out[3806] <= in[514]; 
        out[3807] <= in[1341]; 
        out[3808] <= in[1334]; 
        out[3809] <= in[887]; 
        out[3810] <= in[1258]; 
        out[3811] <= in[3435]; 
        out[3812] <= in[3879]; 
        out[3813] <= in[894]; 
        out[3814] <= in[3247]; 
        out[3815] <= in[2613]; 
        out[3816] <= in[1011]; 
        out[3817] <= in[204]; 
        out[3818] <= in[745]; 
        out[3819] <= in[2159]; 
        out[3820] <= in[2023]; 
        out[3821] <= in[493]; 
        out[3822] <= in[1190]; 
        out[3823] <= in[2110]; 
        out[3824] <= in[3581]; 
        out[3825] <= in[2547]; 
        out[3826] <= in[1310]; 
        out[3827] <= in[457]; 
        out[3828] <= in[2863]; 
        out[3829] <= in[2794]; 
        out[3830] <= in[3295]; 
        out[3831] <= in[409]; 
        out[3832] <= in[1046]; 
        out[3833] <= in[2561]; 
        out[3834] <= in[3413]; 
        out[3835] <= in[4078]; 
        out[3836] <= in[2625]; 
        out[3837] <= in[73]; 
        out[3838] <= in[2282]; 
        out[3839] <= in[139]; 
        out[3840] <= in[2083]; 
        out[3841] <= in[2878]; 
        out[3842] <= in[1145]; 
        out[3843] <= in[2216]; 
        out[3844] <= in[1392]; 
        out[3845] <= in[2207]; 
        out[3846] <= in[3007]; 
        out[3847] <= in[339]; 
        out[3848] <= in[1902]; 
        out[3849] <= in[3593]; 
        out[3850] <= in[1796]; 
        out[3851] <= in[3890]; 
        out[3852] <= in[3461]; 
        out[3853] <= in[2343]; 
        out[3854] <= in[4058]; 
        out[3855] <= in[1186]; 
        out[3856] <= in[1266]; 
        out[3857] <= in[2985]; 
        out[3858] <= in[513]; 
        out[3859] <= in[3537]; 
        out[3860] <= in[3533]; 
        out[3861] <= in[1702]; 
        out[3862] <= in[712]; 
        out[3863] <= in[2767]; 
        out[3864] <= in[2823]; 
        out[3865] <= in[3734]; 
        out[3866] <= in[3659]; 
        out[3867] <= in[2439]; 
        out[3868] <= in[1283]; 
        out[3869] <= in[2093]; 
        out[3870] <= in[1863]; 
        out[3871] <= in[699]; 
        out[3872] <= in[3582]; 
        out[3873] <= in[1518]; 
        out[3874] <= in[1299]; 
        out[3875] <= in[2273]; 
        out[3876] <= in[3130]; 
        out[3877] <= in[1671]; 
        out[3878] <= in[1913]; 
        out[3879] <= in[2495]; 
        out[3880] <= in[594]; 
        out[3881] <= in[1090]; 
        out[3882] <= in[528]; 
        out[3883] <= in[2121]; 
        out[3884] <= in[3699]; 
        out[3885] <= in[666]; 
        out[3886] <= in[411]; 
        out[3887] <= in[2798]; 
        out[3888] <= in[2557]; 
        out[3889] <= in[3637]; 
        out[3890] <= in[2637]; 
        out[3891] <= in[1251]; 
        out[3892] <= in[3658]; 
        out[3893] <= in[1132]; 
        out[3894] <= in[2041]; 
        out[3895] <= in[3984]; 
        out[3896] <= in[1212]; 
        out[3897] <= in[759]; 
        out[3898] <= in[1263]; 
        out[3899] <= in[2697]; 
        out[3900] <= in[929]; 
        out[3901] <= in[3762]; 
        out[3902] <= in[1692]; 
        out[3903] <= in[1899]; 
        out[3904] <= in[1342]; 
        out[3905] <= in[544]; 
        out[3906] <= in[2302]; 
        out[3907] <= in[3680]; 
        out[3908] <= in[848]; 
        out[3909] <= in[3263]; 
        out[3910] <= in[2236]; 
        out[3911] <= in[151]; 
        out[3912] <= in[2317]; 
        out[3913] <= in[266]; 
        out[3914] <= in[1644]; 
        out[3915] <= in[1928]; 
        out[3916] <= in[1386]; 
        out[3917] <= in[1393]; 
        out[3918] <= in[3038]; 
        out[3919] <= in[1757]; 
        out[3920] <= in[3249]; 
        out[3921] <= in[1423]; 
        out[3922] <= in[3379]; 
        out[3923] <= in[2151]; 
        out[3924] <= in[226]; 
        out[3925] <= in[390]; 
        out[3926] <= in[2789]; 
        out[3927] <= in[957]; 
        out[3928] <= in[2936]; 
        out[3929] <= in[172]; 
        out[3930] <= in[2438]; 
        out[3931] <= in[1303]; 
        out[3932] <= in[3516]; 
        out[3933] <= in[2903]; 
        out[3934] <= in[2283]; 
        out[3935] <= in[4013]; 
        out[3936] <= in[1747]; 
        out[3937] <= in[3394]; 
        out[3938] <= in[3875]; 
        out[3939] <= in[2434]; 
        out[3940] <= in[3419]; 
        out[3941] <= in[3793]; 
        out[3942] <= in[1961]; 
        out[3943] <= in[229]; 
        out[3944] <= in[3824]; 
        out[3945] <= in[3982]; 
        out[3946] <= in[2004]; 
        out[3947] <= in[2639]; 
        out[3948] <= in[1804]; 
        out[3949] <= in[944]; 
        out[3950] <= in[869]; 
        out[3951] <= in[3180]; 
        out[3952] <= in[2872]; 
        out[3953] <= in[427]; 
        out[3954] <= in[467]; 
        out[3955] <= in[3331]; 
        out[3956] <= in[37]; 
        out[3957] <= in[338]; 
        out[3958] <= in[3170]; 
        out[3959] <= in[2281]; 
        out[3960] <= in[2653]; 
        out[3961] <= in[1628]; 
        out[3962] <= in[2733]; 
        out[3963] <= in[2735]; 
        out[3964] <= in[3035]; 
        out[3965] <= in[2326]; 
        out[3966] <= in[381]; 
        out[3967] <= in[3311]; 
        out[3968] <= in[1414]; 
        out[3969] <= in[2912]; 
        out[3970] <= in[466]; 
        out[3971] <= in[656]; 
        out[3972] <= in[3724]; 
        out[3973] <= in[2500]; 
        out[3974] <= in[902]; 
        out[3975] <= in[248]; 
        out[3976] <= in[3152]; 
        out[3977] <= in[1442]; 
        out[3978] <= in[3321]; 
        out[3979] <= in[3075]; 
        out[3980] <= in[1214]; 
        out[3981] <= in[2835]; 
        out[3982] <= in[2638]; 
        out[3983] <= in[471]; 
        out[3984] <= in[3725]; 
        out[3985] <= in[3027]; 
        out[3986] <= in[2382]; 
        out[3987] <= in[1802]; 
        out[3988] <= in[3306]; 
        out[3989] <= in[2130]; 
        out[3990] <= in[2967]; 
        out[3991] <= in[3037]; 
        out[3992] <= in[3647]; 
        out[3993] <= in[1219]; 
        out[3994] <= in[4084]; 
        out[3995] <= in[453]; 
        out[3996] <= in[3345]; 
        out[3997] <= in[2415]; 
        out[3998] <= in[2484]; 
        out[3999] <= in[1478]; 
        out[4000] <= in[3962]; 
        out[4001] <= in[3868]; 
        out[4002] <= in[128]; 
        out[4003] <= in[3238]; 
        out[4004] <= in[4070]; 
        out[4005] <= in[3326]; 
        out[4006] <= in[1250]; 
        out[4007] <= in[159]; 
        out[4008] <= in[1381]; 
        out[4009] <= in[237]; 
        out[4010] <= in[305]; 
        out[4011] <= in[2116]; 
        out[4012] <= in[264]; 
        out[4013] <= in[3254]; 
        out[4014] <= in[1216]; 
        out[4015] <= in[1191]; 
        out[4016] <= in[2264]; 
        out[4017] <= in[219]; 
        out[4018] <= in[1551]; 
        out[4019] <= in[1748]; 
        out[4020] <= in[195]; 
        out[4021] <= in[3333]; 
        out[4022] <= in[971]; 
        out[4023] <= in[976]; 
        out[4024] <= in[3036]; 
        out[4025] <= in[3266]; 
        out[4026] <= in[3592]; 
        out[4027] <= in[2719]; 
        out[4028] <= in[3219]; 
        out[4029] <= in[2660]; 
        out[4030] <= in[3960]; 
        out[4031] <= in[2487]; 
        out[4032] <= in[353]; 
        out[4033] <= in[3847]; 
        out[4034] <= in[1549]; 
        out[4035] <= in[3876]; 
        out[4036] <= in[3818]; 
        out[4037] <= in[2015]; 
        out[4038] <= in[2091]; 
        out[4039] <= in[3674]; 
        out[4040] <= in[2440]; 
        out[4041] <= in[1463]; 
        out[4042] <= in[3934]; 
        out[4043] <= in[3656]; 
        out[4044] <= in[2362]; 
        out[4045] <= in[2289]; 
        out[4046] <= in[1468]; 
        out[4047] <= in[2092]; 
        out[4048] <= in[2488]; 
        out[4049] <= in[2319]; 
        out[4050] <= in[3505]; 
        out[4051] <= in[626]; 
        out[4052] <= in[2470]; 
        out[4053] <= in[521]; 
        out[4054] <= in[2467]; 
        out[4055] <= in[2400]; 
        out[4056] <= in[3622]; 
        out[4057] <= in[2480]; 
        out[4058] <= in[2444]; 
        out[4059] <= in[595]; 
        out[4060] <= in[3046]; 
        out[4061] <= in[2056]; 
        out[4062] <= in[1277]; 
        out[4063] <= in[244]; 
        out[4064] <= in[1008]; 
        out[4065] <= in[1473]; 
        out[4066] <= in[212]; 
        out[4067] <= in[3388]; 
        out[4068] <= in[477]; 
        out[4069] <= in[3823]; 
        out[4070] <= in[3517]; 
        out[4071] <= in[3862]; 
        out[4072] <= in[2229]; 
        out[4073] <= in[2721]; 
        out[4074] <= in[2295]; 
        out[4075] <= in[3920]; 
        out[4076] <= in[3790]; 
        out[4077] <= in[1003]; 
        out[4078] <= in[3252]; 
        out[4079] <= in[582]; 
        out[4080] <= in[1517]; 
        out[4081] <= in[1858]; 
        out[4082] <= in[3104]; 
        out[4083] <= in[805]; 
        out[4084] <= in[3682]; 
        out[4085] <= in[3365]; 
        out[4086] <= in[1358]; 
        out[4087] <= in[1709]; 
        out[4088] <= in[625]; 
        out[4089] <= in[834]; 
        out[4090] <= in[2405]; 
        out[4091] <= in[2321]; 
        out[4092] <= in[1821]; 
        out[4093] <= in[3957]; 
        out[4094] <= in[1346]; 
        out[4095] <= in[3837];   
    end

endmodule