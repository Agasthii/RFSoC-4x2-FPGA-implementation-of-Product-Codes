`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/11/2024 05:00:27 PM
// Design Name: 
// Module Name: PC_encoding_block_ebch_256_239
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PC_encoding_block_ebch_256_239 #(
    parameter k = 239,
    parameter n = 256
    )(
    input wire clk,
    input wire reset,
    input wire [4095:0] seed,
    input wire hold_enc,    // Signal from the decoder to start encoding
    output reg store,       // Signal to the datapath to store the encoded codewords in the buffer
    output reg new1,        // Signal to the decoder that a new encoded codeword set is released
    output reg [n-1:0] out_codeword1,
    output reg [n-1:0] out_codeword2,
    output reg [n-1:0] out_codeword3,
    output reg [n-1:0] out_codeword4,
    output reg [n-1:0] out_codeword5,
    output reg [n-1:0] out_codeword6,
    output reg [n-1:0] out_codeword7,
    output reg [n-1:0] out_codeword8,
    output reg [n-1:0] out_codeword9,
    output reg [n-1:0] out_codeword10,
    output reg [n-1:0] out_codeword11,
    output reg [n-1:0] out_codeword12,
    output reg [n-1:0] out_codeword13,
    output reg [n-1:0] out_codeword14,
    output reg [n-1:0] out_codeword15,
    output reg [n-1:0] out_codeword16
    );
    
    // The control variables
    reg [3:0] row_counter = 4'b0; // Counts how many codewords have been stored in the register
    reg [4:0] col_counter = 5'b0; // Counts how many codewords have already given as output
    reg [3:0] set_id = 4'b0;
    reg [1:0] start = 2'b0;
    reg row = 1'b1;
    
    // The outputs from the bit_gen
    wire [k-1:0] bits1;
    wire [k-1:0] bits2;
    wire [k-1:0] bits3;
    wire [k-1:0] bits4;
    wire [k-1:0] bits5;
    wire [k-1:0] bits6;
    wire [k-1:0] bits7;
    wire [k-1:0] bits8;
    wire [k-1:0] bits9;
    wire [k-1:0] bits10;
    wire [k-1:0] bits11;
    wire [k-1:0] bits12;
    wire [k-1:0] bits13;
    wire [k-1:0] bits14;
    wire [k-1:0] bits15;
    wire [k-1:0] bits16;
    
    // The inputs to the encoders
    reg [k-1:0] in_bits1;
    reg [k-1:0] in_bits2;
    reg [k-1:0] in_bits3;
    reg [k-1:0] in_bits4;
    reg [k-1:0] in_bits5;
    reg [k-1:0] in_bits6;
    reg [k-1:0] in_bits7;
    reg [k-1:0] in_bits8;
    reg [k-1:0] in_bits9;
    reg [k-1:0] in_bits10;
    reg [k-1:0] in_bits11;
    reg [k-1:0] in_bits12;
    reg [k-1:0] in_bits13;
    reg [k-1:0] in_bits14;
    reg [k-1:0] in_bits15;
    reg [k-1:0] in_bits16;
    
    // The buffer to store the outputs from the row encoding
    reg [n*15-1:0] codeword_reg1;
    reg [n*15-1:0] codeword_reg2;
    reg [n*15-1:0] codeword_reg3;
    reg [n*15-1:0] codeword_reg4;
    reg [n*15-1:0] codeword_reg5;
    reg [n*15-1:0] codeword_reg6;
    reg [n*15-1:0] codeword_reg7;
    reg [n*15-1:0] codeword_reg8;
    reg [n*15-1:0] codeword_reg9;
    reg [n*15-1:0] codeword_reg10;
    reg [n*15-1:0] codeword_reg11;
    reg [n*15-1:0] codeword_reg12;
    reg [n*15-1:0] codeword_reg13;
    reg [n*15-1:0] codeword_reg14;
    reg [n*15-1:0] codeword_reg15;
    reg [n*15-1:0] codeword_reg16;  
    
    // The outputs from the row encoding
    wire [n-1:0] codeword1;
    wire [n-1:0] codeword2;
    wire [n-1:0] codeword3;
    wire [n-1:0] codeword4;
    wire [n-1:0] codeword5;
    wire [n-1:0] codeword6;
    wire [n-1:0] codeword7;
    wire [n-1:0] codeword8;
    wire [n-1:0] codeword9;
    wire [n-1:0] codeword10;
    wire [n-1:0] codeword11;
    wire [n-1:0] codeword12;
    wire [n-1:0] codeword13;
    wire [n-1:0] codeword14;
    wire [n-1:0] codeword15;
    wire [n-1:0] codeword16;
    
    bit_gen_PC bit_gen(
        .clk(clk),
        .reset(reset),
        .seed(seed),
        .bits1(bits1),
        .bits2(bits2),
        .bits3(bits3),
        .bits4(bits4),
        .bits5(bits5),
        .bits6(bits6),
        .bits7(bits7),
        .bits8(bits8),
        .bits9(bits9),
        .bits10(bits10),
        .bits11(bits11),
        .bits12(bits12),
        .bits13(bits13),
        .bits14(bits14),
        .bits15(bits15),
        .bits16(bits16)
        );
          
    
    bchencoder_256_239_PC encoder(
        .clk(clk),
        .reset(reset),
        .bits1(in_bits1),
        .bits2(in_bits2),
        .bits3(in_bits3),
        .bits4(in_bits4),
        .bits5(in_bits5),
        .bits6(in_bits6),
        .bits7(in_bits7),
        .bits8(in_bits8),
        .bits9(in_bits9),
        .bits10(in_bits10),
        .bits11(in_bits11),
        .bits12(in_bits12),
        .bits13(in_bits13),
        .bits14(in_bits14),
        .bits15(in_bits15),
        .bits16(in_bits16),
        .codeword1(codeword1),
        .codeword2(codeword2),
        .codeword3(codeword3),
        .codeword4(codeword4),
        .codeword5(codeword5),
        .codeword6(codeword6),
        .codeword7(codeword7),
        .codeword8(codeword8),
        .codeword9(codeword9),
        .codeword10(codeword10),
        .codeword11(codeword11),
        .codeword12(codeword12),
        .codeword13(codeword13),
        .codeword14(codeword14),
        .codeword15(codeword15),
        .codeword16(codeword16)
    );
    
    always@(posedge clk) begin
        // If the system is OFF
        if (!reset) begin
            row_counter <= 4'b0;
            col_counter <= 5'b0;
            set_id <= 4'b0;
            start <= 2'b0;
            new1 <= 1'b0;
            
        // If the system is ON
        end else begin
        
            //// Start of the encoding ////
            if (hold_enc) begin
            
                // if the encoding is allowed from the decoder
                if (start == 2'b11) begin
                
                    //// Start of the row encoding ////
                    if (row == 1'b1) begin
                    
                        // If the row encoding is for the first 14
                        if (row_counter < 4'd14) begin        
                            
                            // Give the generated bits to the row encoder
                            in_bits1  <= bits1;
                            in_bits2  <= bits2;
                            in_bits3  <= bits3;
                            in_bits4  <= bits4;
                            in_bits5  <= bits5;
                            in_bits6  <= bits6;
                            in_bits7  <= bits7;
                            in_bits8  <= bits8;
                            in_bits9  <= bits9;
                            in_bits10 <= bits10;
                            in_bits11 <= bits11;
                            in_bits12 <= bits12;
                            in_bits13 <= bits13;
                            in_bits14 <= bits14;
                            in_bits15 <= bits15;
                            in_bits16 <= bits16;
                            
                            // Shift the buffer to store the row encoded codewords
                            codeword_reg1[(set_id)*n  +: n] <= codeword1;
                            codeword_reg2[(set_id)*n  +: n] <= codeword2;
                            codeword_reg3[(set_id)*n  +: n] <= codeword3;
                            codeword_reg4[(set_id)*n  +: n] <= codeword4;
                            codeword_reg5[(set_id)*n  +: n] <= codeword5;
                            codeword_reg6[(set_id)*n  +: n] <= codeword6;
                            codeword_reg7[(set_id)*n  +: n] <= codeword7;
                            codeword_reg8[(set_id)*n  +: n] <= codeword8;
                            codeword_reg9[(set_id)*n  +: n] <= codeword9;
                            codeword_reg10[(set_id)*n +: n] <= codeword10;
                            codeword_reg11[(set_id)*n +: n] <= codeword11;
                            codeword_reg12[(set_id)*n +: n] <= codeword12;
                            codeword_reg13[(set_id)*n +: n] <= codeword13;
                            codeword_reg14[(set_id)*n +: n] <= codeword14;
                            codeword_reg15[(set_id)*n +: n] <= codeword15;
                            codeword_reg16[(set_id)*n +: n] <= codeword16;
                            
                            // Output x as the encoded codewords
                            out_codeword1  <= 'bx;
                            out_codeword2  <= 'bx;
                            out_codeword3  <= 'bx;
                            out_codeword4  <= 'bx;
                            out_codeword5  <= 'bx;
                            out_codeword6  <= 'bx;
                            out_codeword7  <= 'bx;
                            out_codeword8  <= 'bx;
                            out_codeword9  <= 'bx;
                            out_codeword10 <= 'bx;
                            out_codeword11 <= 'bx;
                            out_codeword12 <= 'bx;
                            out_codeword13 <= 'bx;
                            out_codeword14 <= 'bx;
                            out_codeword15 <= 'bx;
                            out_codeword16 <= 'bx;
                            
                            // Update the control variables
                            set_id <= set_id + 4'b1;
                            row_counter <= row_counter + 1;
                            new1 <= 1'b0;
                            store <= 1'b0;
                        
                        // If the row encoding is for the 15th codeword                 
                        end else begin 
                            
//                            in_bits1  <= {codeword16[0], codeword15[0], codeword14[0], codeword13[0], codeword12[0], codeword11[0], codeword10[0], codeword9[0], codeword8[0], codeword7[0], codeword6[0], codeword5[0], codeword4[0], codeword3[0], codeword2[0], codeword1[0], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits2  <= {codeword16[1], codeword15[1], codeword14[1], codeword13[1], codeword12[1], codeword11[1], codeword10[1], codeword9[1], codeword8[1], codeword7[1], codeword6[1], codeword5[1], codeword4[1], codeword3[1], codeword2[1], codeword1[1], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits3  <= {codeword16[2], codeword15[2], codeword14[2], codeword13[2], codeword12[2], codeword11[2], codeword10[2], codeword9[2], codeword8[2], codeword7[2], codeword6[2], codeword5[2], codeword4[2], codeword3[2], codeword2[2], codeword1[2], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits4  <= {codeword16[3], codeword15[3], codeword14[3], codeword13[3], codeword12[3], codeword11[3], codeword10[3], codeword9[3], codeword8[3], codeword7[3], codeword6[3], codeword5[3], codeword4[3], codeword3[3], codeword2[3], codeword1[3], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits5  <= {codeword16[4], codeword15[4], codeword14[4], codeword13[4], codeword12[4], codeword11[4], codeword10[4], codeword9[4], codeword8[4], codeword7[4], codeword6[4], codeword5[4], codeword4[4], codeword3[4], codeword2[4], codeword1[4], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits6  <= {codeword16[5], codeword15[5], codeword14[5], codeword13[5], codeword12[5], codeword11[5], codeword10[5], codeword9[5], codeword8[5], codeword7[5], codeword6[5], codeword5[5], codeword4[5], codeword3[5], codeword2[5], codeword1[5], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits7  <= {codeword16[6], codeword15[6], codeword14[6], codeword13[6], codeword12[6], codeword11[6], codeword10[6], codeword9[6], codeword8[6], codeword7[6], codeword6[6], codeword5[6], codeword4[6], codeword3[6], codeword2[6], codeword1[6], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits8  <= {codeword16[7], codeword15[7], codeword14[7], codeword13[7], codeword12[7], codeword11[7], codeword10[7], codeword9[7], codeword8[7], codeword7[7], codeword6[7], codeword5[7], codeword4[7], codeword3[7], codeword2[7], codeword1[7], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits9  <= {codeword16[8], codeword15[8], codeword14[8], codeword13[8], codeword12[8], codeword11[8], codeword10[8], codeword9[8], codeword8[8], codeword7[8], codeword6[8], codeword5[8], codeword4[8], codeword3[8], codeword2[8], codeword1[8], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits10 <= {codeword16[9], codeword15[9], codeword14[9], codeword13[9], codeword12[9], codeword11[9], codeword10[9], codeword9[9], codeword8[9], codeword7[9], codeword6[9], codeword5[9], codeword4[9], codeword3[9], codeword2[9], codeword1[9], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits11 <= {codeword16[10], codeword15[10], codeword14[10], codeword13[10], codeword12[10], codeword11[10], codeword10[10], codeword9[10], codeword8[10], codeword7[10], codeword6[10], codeword5[10], codeword4[10], codeword3[10], codeword2[10], codeword1[10], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits12 <= {codeword16[11], codeword15[11], codeword14[11], codeword13[11], codeword12[11], codeword11[11], codeword10[11], codeword9[11], codeword8[11], codeword7[11], codeword6[11], codeword5[11], codeword4[11], codeword3[11], codeword2[11], codeword1[11], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits13 <= {codeword16[12], codeword15[12], codeword14[12], codeword13[12], codeword12[12], codeword11[12], codeword10[12], codeword9[12], codeword8[12], codeword7[12], codeword6[12], codeword5[12], codeword4[12], codeword3[12], codeword2[12], codeword1[12], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits14 <= {codeword16[13], codeword15[13], codeword14[13], codeword13[13], codeword12[13], codeword11[13], codeword10[13], codeword9[13], codeword8[13], codeword7[13], codeword6[13], codeword5[13], codeword4[13], codeword3[13], codeword2[13], codeword1[13], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits15 <= {codeword16[14], codeword15[14], codeword14[14], codeword13[14], codeword12[14], codeword11[14], codeword10[14], codeword9[14], codeword8[14], codeword7[14], codeword6[14], codeword5[14], codeword4[14], codeword3[14], codeword2[14], codeword1[14], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
//                            in_bits16 <= {codeword16[15], codeword15[15], codeword14[15], codeword13[15], codeword12[15], codeword11[15], codeword10[15], codeword9[15], codeword8[15], codeword7[15], codeword6[15], codeword5[15], codeword4[15], codeword3[15], codeword2[15], codeword1[15], codeword_reg16[256*13], codeword_reg15[256*13], codeword_reg14[256*13], codeword_reg13[256*13], codeword_reg12[256*13], codeword_reg11[256*13], codeword_reg10[256*13], codeword_reg9[256*13], codeword_reg8[256*13], codeword_reg7[256*13], codeword_reg6[256*13], codeword_reg5[256*13], codeword_reg4[256*13], codeword_reg3[256*13], codeword_reg2[256*13], codeword_reg1[256*13], codeword_reg16[256*12], codeword_reg15[256*12], codeword_reg14[256*12], codeword_reg13[256*12], codeword_reg12[256*12], codeword_reg11[256*12], codeword_reg10[256*12], codeword_reg9[256*12], codeword_reg8[256*12], codeword_reg7[256*12], codeword_reg6[256*12], codeword_reg5[256*12], codeword_reg4[256*12], codeword_reg3[256*12], codeword_reg2[256*12], codeword_reg1[256*12], codeword_reg16[256*11], codeword_reg15[256*11], codeword_reg14[256*11], codeword_reg13[256*11], codeword_reg12[256*11], codeword_reg11[256*11], codeword_reg10[256*11], codeword_reg9[256*11], codeword_reg8[256*11], codeword_reg7[256*11], codeword_reg6[256*11], codeword_reg5[256*11], codeword_reg4[256*11], codeword_reg3[256*11], codeword_reg2[256*11], codeword_reg1[256*11], codeword_reg16[256*10], codeword_reg15[256*10], codeword_reg14[256*10], codeword_reg13[256*10], codeword_reg12[256*10], codeword_reg11[256*10], codeword_reg10[256*10], codeword_reg9[256*10], codeword_reg8[256*10], codeword_reg7[256*10], codeword_reg6[256*10], codeword_reg5[256*10], codeword_reg4[256*10], codeword_reg3[256*10], codeword_reg2[256*10], codeword_reg1[256*10], codeword_reg16[256*9], codeword_reg15[256*9], codeword_reg14[256*9], codeword_reg13[256*9], codeword_reg12[256*9], codeword_reg11[256*9], codeword_reg10[256*9], codeword_reg9[256*9], codeword_reg8[256*9], codeword_reg7[256*9], codeword_reg6[256*9], codeword_reg5[256*9], codeword_reg4[256*9], codeword_reg3[256*9], codeword_reg2[256*9], codeword_reg1[256*9], codeword_reg16[256*8], codeword_reg15[256*8], codeword_reg14[256*8], codeword_reg13[256*8], codeword_reg12[256*8], codeword_reg11[256*8], codeword_reg10[256*8], codeword_reg9[256*8], codeword_reg8[256*8], codeword_reg7[256*8], codeword_reg6[256*8], codeword_reg5[256*8], codeword_reg4[256*8], codeword_reg3[256*8], codeword_reg2[256*8], codeword_reg1[256*8], codeword_reg16[256*7], codeword_reg15[256*7], codeword_reg14[256*7], codeword_reg13[256*7], codeword_reg12[256*7], codeword_reg11[256*7], codeword_reg10[256*7], codeword_reg9[256*7], codeword_reg8[256*7], codeword_reg7[256*7], codeword_reg6[256*7], codeword_reg5[256*7], codeword_reg4[256*7], codeword_reg3[256*7], codeword_reg2[256*7], codeword_reg1[256*7], codeword_reg16[256*6], codeword_reg15[256*6], codeword_reg14[256*6], codeword_reg13[256*6], codeword_reg12[256*6], codeword_reg11[256*6], codeword_reg10[256*6], codeword_reg9[256*6], codeword_reg8[256*6], codeword_reg7[256*6], codeword_reg6[256*6], codeword_reg5[256*6], codeword_reg4[256*6], codeword_reg3[256*6], codeword_reg2[256*6], codeword_reg1[256*6], codeword_reg16[256*5], codeword_reg15[256*5], codeword_reg14[256*5], codeword_reg13[256*5], codeword_reg12[256*5], codeword_reg11[256*5], codeword_reg10[256*5], codeword_reg9[256*5], codeword_reg8[256*5], codeword_reg7[256*5], codeword_reg6[256*5], codeword_reg5[256*5], codeword_reg4[256*5], codeword_reg3[256*5], codeword_reg2[256*5], codeword_reg1[256*5], codeword_reg16[256*4], codeword_reg15[256*4], codeword_reg14[256*4], codeword_reg13[256*4], codeword_reg12[256*4], codeword_reg11[256*4], codeword_reg10[256*4], codeword_reg9[256*4], codeword_reg8[256*4], codeword_reg7[256*4], codeword_reg6[256*4], codeword_reg5[256*4], codeword_reg4[256*4], codeword_reg3[256*4], codeword_reg2[256*4], codeword_reg1[256*4], codeword_reg16[256*3], codeword_reg15[256*3], codeword_reg14[256*3], codeword_reg13[256*3], codeword_reg12[256*3], codeword_reg11[256*3], codeword_reg10[256*3], codeword_reg9[256*3], codeword_reg8[256*3], codeword_reg7[256*3], codeword_reg6[256*3], codeword_reg5[256*3], codeword_reg4[256*3], codeword_reg3[256*3], codeword_reg2[256*3], codeword_reg1[256*3], codeword_reg16[256*2], codeword_reg15[256*2], codeword_reg14[256*2], codeword_reg13[256*2], codeword_reg12[256*2], codeword_reg11[256*2], codeword_reg10[256*2], codeword_reg9[256*2], codeword_reg8[256*2], codeword_reg7[256*2], codeword_reg6[256*2], codeword_reg5[256*2], codeword_reg4[256*2], codeword_reg3[256*2], codeword_reg2[256*2], codeword_reg1[256*2], codeword_reg16[256*1], codeword_reg15[256*1], codeword_reg14[256*1], codeword_reg13[256*1], codeword_reg12[256*1], codeword_reg11[256*1], codeword_reg10[256*1], codeword_reg9[256*1], codeword_reg8[256*1], codeword_reg7[256*1], codeword_reg6[256*1], codeword_reg5[256*1], codeword_reg4[256*1], codeword_reg3[256*1], codeword_reg2[256*1], codeword_reg1[256*1], codeword_reg16[256*0], codeword_reg15[256*0], codeword_reg14[256*0], codeword_reg13[256*0], codeword_reg12[256*0], codeword_reg11[256*0], codeword_reg10[256*0], codeword_reg9[256*0], codeword_reg8[256*0], codeword_reg7[256*0], codeword_reg6[256*0], codeword_reg5[256*0], codeword_reg4[256*0], codeword_reg3[256*0], codeword_reg2[256*0], codeword_reg1[256*0]};
                            
                            in_bits1 <= {codeword16[0], codeword15[0], codeword14[0], codeword13[0], codeword12[0], codeword11[0], codeword10[0], codeword9[0], codeword8[0], codeword7[0], codeword6[0], codeword5[0], codeword4[0], codeword3[0], codeword2[0], codeword1[0], codeword_reg16[256*13+0], codeword_reg15[256*13+0], codeword_reg14[256*13+0], codeword_reg13[256*13+0], codeword_reg12[256*13+0], codeword_reg11[256*13+0], codeword_reg10[256*13+0], codeword_reg9[256*13+0], codeword_reg8[256*13+0], codeword_reg7[256*13+0], codeword_reg6[256*13+0], codeword_reg5[256*13+0], codeword_reg4[256*13+0], codeword_reg3[256*13+0], codeword_reg2[256*13+0], codeword_reg1[256*13+0], codeword_reg16[256*12+0], codeword_reg15[256*12+0], codeword_reg14[256*12+0], codeword_reg13[256*12+0], codeword_reg12[256*12+0], codeword_reg11[256*12+0], codeword_reg10[256*12+0], codeword_reg9[256*12+0], codeword_reg8[256*12+0], codeword_reg7[256*12+0], codeword_reg6[256*12+0], codeword_reg5[256*12+0], codeword_reg4[256*12+0], codeword_reg3[256*12+0], codeword_reg2[256*12+0], codeword_reg1[256*12+0], codeword_reg16[256*11+0], codeword_reg15[256*11+0], codeword_reg14[256*11+0], codeword_reg13[256*11+0], codeword_reg12[256*11+0], codeword_reg11[256*11+0], codeword_reg10[256*11+0], codeword_reg9[256*11+0], codeword_reg8[256*11+0], codeword_reg7[256*11+0], codeword_reg6[256*11+0], codeword_reg5[256*11+0], codeword_reg4[256*11+0], codeword_reg3[256*11+0], codeword_reg2[256*11+0], codeword_reg1[256*11+0], codeword_reg16[256*10+0], codeword_reg15[256*10+0], codeword_reg14[256*10+0], codeword_reg13[256*10+0], codeword_reg12[256*10+0], codeword_reg11[256*10+0], codeword_reg10[256*10+0], codeword_reg9[256*10+0], codeword_reg8[256*10+0], codeword_reg7[256*10+0], codeword_reg6[256*10+0], codeword_reg5[256*10+0], codeword_reg4[256*10+0], codeword_reg3[256*10+0], codeword_reg2[256*10+0], codeword_reg1[256*10+0], codeword_reg16[256*9+0], codeword_reg15[256*9+0], codeword_reg14[256*9+0], codeword_reg13[256*9+0], codeword_reg12[256*9+0], codeword_reg11[256*9+0], codeword_reg10[256*9+0], codeword_reg9[256*9+0], codeword_reg8[256*9+0], codeword_reg7[256*9+0], codeword_reg6[256*9+0], codeword_reg5[256*9+0], codeword_reg4[256*9+0], codeword_reg3[256*9+0], codeword_reg2[256*9+0], codeword_reg1[256*9+0], codeword_reg16[256*8+0], codeword_reg15[256*8+0], codeword_reg14[256*8+0], codeword_reg13[256*8+0], codeword_reg12[256*8+0], codeword_reg11[256*8+0], codeword_reg10[256*8+0], codeword_reg9[256*8+0], codeword_reg8[256*8+0], codeword_reg7[256*8+0], codeword_reg6[256*8+0], codeword_reg5[256*8+0], codeword_reg4[256*8+0], codeword_reg3[256*8+0], codeword_reg2[256*8+0], codeword_reg1[256*8+0], codeword_reg16[256*7+0], codeword_reg15[256*7+0], codeword_reg14[256*7+0], codeword_reg13[256*7+0], codeword_reg12[256*7+0], codeword_reg11[256*7+0], codeword_reg10[256*7+0], codeword_reg9[256*7+0], codeword_reg8[256*7+0], codeword_reg7[256*7+0], codeword_reg6[256*7+0], codeword_reg5[256*7+0], codeword_reg4[256*7+0], codeword_reg3[256*7+0], codeword_reg2[256*7+0], codeword_reg1[256*7+0], codeword_reg16[256*6+0], codeword_reg15[256*6+0], codeword_reg14[256*6+0], codeword_reg13[256*6+0], codeword_reg12[256*6+0], codeword_reg11[256*6+0], codeword_reg10[256*6+0], codeword_reg9[256*6+0], codeword_reg8[256*6+0], codeword_reg7[256*6+0], codeword_reg6[256*6+0], codeword_reg5[256*6+0], codeword_reg4[256*6+0], codeword_reg3[256*6+0], codeword_reg2[256*6+0], codeword_reg1[256*6+0], codeword_reg16[256*5+0], codeword_reg15[256*5+0], codeword_reg14[256*5+0], codeword_reg13[256*5+0], codeword_reg12[256*5+0], codeword_reg11[256*5+0], codeword_reg10[256*5+0], codeword_reg9[256*5+0], codeword_reg8[256*5+0], codeword_reg7[256*5+0], codeword_reg6[256*5+0], codeword_reg5[256*5+0], codeword_reg4[256*5+0], codeword_reg3[256*5+0], codeword_reg2[256*5+0], codeword_reg1[256*5+0], codeword_reg16[256*4+0], codeword_reg15[256*4+0], codeword_reg14[256*4+0], codeword_reg13[256*4+0], codeword_reg12[256*4+0], codeword_reg11[256*4+0], codeword_reg10[256*4+0], codeword_reg9[256*4+0], codeword_reg8[256*4+0], codeword_reg7[256*4+0], codeword_reg6[256*4+0], codeword_reg5[256*4+0], codeword_reg4[256*4+0], codeword_reg3[256*4+0], codeword_reg2[256*4+0], codeword_reg1[256*4+0], codeword_reg16[256*3+0], codeword_reg15[256*3+0], codeword_reg14[256*3+0], codeword_reg13[256*3+0], codeword_reg12[256*3+0], codeword_reg11[256*3+0], codeword_reg10[256*3+0], codeword_reg9[256*3+0], codeword_reg8[256*3+0], codeword_reg7[256*3+0], codeword_reg6[256*3+0], codeword_reg5[256*3+0], codeword_reg4[256*3+0], codeword_reg3[256*3+0], codeword_reg2[256*3+0], codeword_reg1[256*3+0], codeword_reg16[256*2+0], codeword_reg15[256*2+0], codeword_reg14[256*2+0], codeword_reg13[256*2+0], codeword_reg12[256*2+0], codeword_reg11[256*2+0], codeword_reg10[256*2+0], codeword_reg9[256*2+0], codeword_reg8[256*2+0], codeword_reg7[256*2+0], codeword_reg6[256*2+0], codeword_reg5[256*2+0], codeword_reg4[256*2+0], codeword_reg3[256*2+0], codeword_reg2[256*2+0], codeword_reg1[256*2+0], codeword_reg16[256*1+0], codeword_reg15[256*1+0], codeword_reg14[256*1+0], codeword_reg13[256*1+0], codeword_reg12[256*1+0], codeword_reg11[256*1+0], codeword_reg10[256*1+0], codeword_reg9[256*1+0], codeword_reg8[256*1+0], codeword_reg7[256*1+0], codeword_reg6[256*1+0], codeword_reg5[256*1+0], codeword_reg4[256*1+0], codeword_reg3[256*1+0], codeword_reg2[256*1+0], codeword_reg1[256*1+0], codeword_reg16[256*0+0], codeword_reg15[256*0+0], codeword_reg14[256*0+0], codeword_reg13[256*0+0], codeword_reg12[256*0+0], codeword_reg11[256*0+0], codeword_reg10[256*0+0], codeword_reg9[256*0+0], codeword_reg8[256*0+0], codeword_reg7[256*0+0], codeword_reg6[256*0+0], codeword_reg5[256*0+0], codeword_reg4[256*0+0], codeword_reg3[256*0+0], codeword_reg2[256*0+0], codeword_reg1[256*0+0]};
                                in_bits2 <= {codeword16[1], codeword15[1], codeword14[1], codeword13[1], codeword12[1], codeword11[1], codeword10[1], codeword9[1], codeword8[1], codeword7[1], codeword6[1], codeword5[1], codeword4[1], codeword3[1], codeword2[1], codeword1[1], codeword_reg16[256*13+1], codeword_reg15[256*13+1], codeword_reg14[256*13+1], codeword_reg13[256*13+1], codeword_reg12[256*13+1], codeword_reg11[256*13+1], codeword_reg10[256*13+1], codeword_reg9[256*13+1], codeword_reg8[256*13+1], codeword_reg7[256*13+1], codeword_reg6[256*13+1], codeword_reg5[256*13+1], codeword_reg4[256*13+1], codeword_reg3[256*13+1], codeword_reg2[256*13+1], codeword_reg1[256*13+1], codeword_reg16[256*12+1], codeword_reg15[256*12+1], codeword_reg14[256*12+1], codeword_reg13[256*12+1], codeword_reg12[256*12+1], codeword_reg11[256*12+1], codeword_reg10[256*12+1], codeword_reg9[256*12+1], codeword_reg8[256*12+1], codeword_reg7[256*12+1], codeword_reg6[256*12+1], codeword_reg5[256*12+1], codeword_reg4[256*12+1], codeword_reg3[256*12+1], codeword_reg2[256*12+1], codeword_reg1[256*12+1], codeword_reg16[256*11+1], codeword_reg15[256*11+1], codeword_reg14[256*11+1], codeword_reg13[256*11+1], codeword_reg12[256*11+1], codeword_reg11[256*11+1], codeword_reg10[256*11+1], codeword_reg9[256*11+1], codeword_reg8[256*11+1], codeword_reg7[256*11+1], codeword_reg6[256*11+1], codeword_reg5[256*11+1], codeword_reg4[256*11+1], codeword_reg3[256*11+1], codeword_reg2[256*11+1], codeword_reg1[256*11+1], codeword_reg16[256*10+1], codeword_reg15[256*10+1], codeword_reg14[256*10+1], codeword_reg13[256*10+1], codeword_reg12[256*10+1], codeword_reg11[256*10+1], codeword_reg10[256*10+1], codeword_reg9[256*10+1], codeword_reg8[256*10+1], codeword_reg7[256*10+1], codeword_reg6[256*10+1], codeword_reg5[256*10+1], codeword_reg4[256*10+1], codeword_reg3[256*10+1], codeword_reg2[256*10+1], codeword_reg1[256*10+1], codeword_reg16[256*9+1], codeword_reg15[256*9+1], codeword_reg14[256*9+1], codeword_reg13[256*9+1], codeword_reg12[256*9+1], codeword_reg11[256*9+1], codeword_reg10[256*9+1], codeword_reg9[256*9+1], codeword_reg8[256*9+1], codeword_reg7[256*9+1], codeword_reg6[256*9+1], codeword_reg5[256*9+1], codeword_reg4[256*9+1], codeword_reg3[256*9+1], codeword_reg2[256*9+1], codeword_reg1[256*9+1], codeword_reg16[256*8+1], codeword_reg15[256*8+1], codeword_reg14[256*8+1], codeword_reg13[256*8+1], codeword_reg12[256*8+1], codeword_reg11[256*8+1], codeword_reg10[256*8+1], codeword_reg9[256*8+1], codeword_reg8[256*8+1], codeword_reg7[256*8+1], codeword_reg6[256*8+1], codeword_reg5[256*8+1], codeword_reg4[256*8+1], codeword_reg3[256*8+1], codeword_reg2[256*8+1], codeword_reg1[256*8+1], codeword_reg16[256*7+1], codeword_reg15[256*7+1], codeword_reg14[256*7+1], codeword_reg13[256*7+1], codeword_reg12[256*7+1], codeword_reg11[256*7+1], codeword_reg10[256*7+1], codeword_reg9[256*7+1], codeword_reg8[256*7+1], codeword_reg7[256*7+1], codeword_reg6[256*7+1], codeword_reg5[256*7+1], codeword_reg4[256*7+1], codeword_reg3[256*7+1], codeword_reg2[256*7+1], codeword_reg1[256*7+1], codeword_reg16[256*6+1], codeword_reg15[256*6+1], codeword_reg14[256*6+1], codeword_reg13[256*6+1], codeword_reg12[256*6+1], codeword_reg11[256*6+1], codeword_reg10[256*6+1], codeword_reg9[256*6+1], codeword_reg8[256*6+1], codeword_reg7[256*6+1], codeword_reg6[256*6+1], codeword_reg5[256*6+1], codeword_reg4[256*6+1], codeword_reg3[256*6+1], codeword_reg2[256*6+1], codeword_reg1[256*6+1], codeword_reg16[256*5+1], codeword_reg15[256*5+1], codeword_reg14[256*5+1], codeword_reg13[256*5+1], codeword_reg12[256*5+1], codeword_reg11[256*5+1], codeword_reg10[256*5+1], codeword_reg9[256*5+1], codeword_reg8[256*5+1], codeword_reg7[256*5+1], codeword_reg6[256*5+1], codeword_reg5[256*5+1], codeword_reg4[256*5+1], codeword_reg3[256*5+1], codeword_reg2[256*5+1], codeword_reg1[256*5+1], codeword_reg16[256*4+1], codeword_reg15[256*4+1], codeword_reg14[256*4+1], codeword_reg13[256*4+1], codeword_reg12[256*4+1], codeword_reg11[256*4+1], codeword_reg10[256*4+1], codeword_reg9[256*4+1], codeword_reg8[256*4+1], codeword_reg7[256*4+1], codeword_reg6[256*4+1], codeword_reg5[256*4+1], codeword_reg4[256*4+1], codeword_reg3[256*4+1], codeword_reg2[256*4+1], codeword_reg1[256*4+1], codeword_reg16[256*3+1], codeword_reg15[256*3+1], codeword_reg14[256*3+1], codeword_reg13[256*3+1], codeword_reg12[256*3+1], codeword_reg11[256*3+1], codeword_reg10[256*3+1], codeword_reg9[256*3+1], codeword_reg8[256*3+1], codeword_reg7[256*3+1], codeword_reg6[256*3+1], codeword_reg5[256*3+1], codeword_reg4[256*3+1], codeword_reg3[256*3+1], codeword_reg2[256*3+1], codeword_reg1[256*3+1], codeword_reg16[256*2+1], codeword_reg15[256*2+1], codeword_reg14[256*2+1], codeword_reg13[256*2+1], codeword_reg12[256*2+1], codeword_reg11[256*2+1], codeword_reg10[256*2+1], codeword_reg9[256*2+1], codeword_reg8[256*2+1], codeword_reg7[256*2+1], codeword_reg6[256*2+1], codeword_reg5[256*2+1], codeword_reg4[256*2+1], codeword_reg3[256*2+1], codeword_reg2[256*2+1], codeword_reg1[256*2+1], codeword_reg16[256*1+1], codeword_reg15[256*1+1], codeword_reg14[256*1+1], codeword_reg13[256*1+1], codeword_reg12[256*1+1], codeword_reg11[256*1+1], codeword_reg10[256*1+1], codeword_reg9[256*1+1], codeword_reg8[256*1+1], codeword_reg7[256*1+1], codeword_reg6[256*1+1], codeword_reg5[256*1+1], codeword_reg4[256*1+1], codeword_reg3[256*1+1], codeword_reg2[256*1+1], codeword_reg1[256*1+1], codeword_reg16[256*0+1], codeword_reg15[256*0+1], codeword_reg14[256*0+1], codeword_reg13[256*0+1], codeword_reg12[256*0+1], codeword_reg11[256*0+1], codeword_reg10[256*0+1], codeword_reg9[256*0+1], codeword_reg8[256*0+1], codeword_reg7[256*0+1], codeword_reg6[256*0+1], codeword_reg5[256*0+1], codeword_reg4[256*0+1], codeword_reg3[256*0+1], codeword_reg2[256*0+1], codeword_reg1[256*0+1]};
                                in_bits3 <= {codeword16[2], codeword15[2], codeword14[2], codeword13[2], codeword12[2], codeword11[2], codeword10[2], codeword9[2], codeword8[2], codeword7[2], codeword6[2], codeword5[2], codeword4[2], codeword3[2], codeword2[2], codeword1[2], codeword_reg16[256*13+2], codeword_reg15[256*13+2], codeword_reg14[256*13+2], codeword_reg13[256*13+2], codeword_reg12[256*13+2], codeword_reg11[256*13+2], codeword_reg10[256*13+2], codeword_reg9[256*13+2], codeword_reg8[256*13+2], codeword_reg7[256*13+2], codeword_reg6[256*13+2], codeword_reg5[256*13+2], codeword_reg4[256*13+2], codeword_reg3[256*13+2], codeword_reg2[256*13+2], codeword_reg1[256*13+2], codeword_reg16[256*12+2], codeword_reg15[256*12+2], codeword_reg14[256*12+2], codeword_reg13[256*12+2], codeword_reg12[256*12+2], codeword_reg11[256*12+2], codeword_reg10[256*12+2], codeword_reg9[256*12+2], codeword_reg8[256*12+2], codeword_reg7[256*12+2], codeword_reg6[256*12+2], codeword_reg5[256*12+2], codeword_reg4[256*12+2], codeword_reg3[256*12+2], codeword_reg2[256*12+2], codeword_reg1[256*12+2], codeword_reg16[256*11+2], codeword_reg15[256*11+2], codeword_reg14[256*11+2], codeword_reg13[256*11+2], codeword_reg12[256*11+2], codeword_reg11[256*11+2], codeword_reg10[256*11+2], codeword_reg9[256*11+2], codeword_reg8[256*11+2], codeword_reg7[256*11+2], codeword_reg6[256*11+2], codeword_reg5[256*11+2], codeword_reg4[256*11+2], codeword_reg3[256*11+2], codeword_reg2[256*11+2], codeword_reg1[256*11+2], codeword_reg16[256*10+2], codeword_reg15[256*10+2], codeword_reg14[256*10+2], codeword_reg13[256*10+2], codeword_reg12[256*10+2], codeword_reg11[256*10+2], codeword_reg10[256*10+2], codeword_reg9[256*10+2], codeword_reg8[256*10+2], codeword_reg7[256*10+2], codeword_reg6[256*10+2], codeword_reg5[256*10+2], codeword_reg4[256*10+2], codeword_reg3[256*10+2], codeword_reg2[256*10+2], codeword_reg1[256*10+2], codeword_reg16[256*9+2], codeword_reg15[256*9+2], codeword_reg14[256*9+2], codeword_reg13[256*9+2], codeword_reg12[256*9+2], codeword_reg11[256*9+2], codeword_reg10[256*9+2], codeword_reg9[256*9+2], codeword_reg8[256*9+2], codeword_reg7[256*9+2], codeword_reg6[256*9+2], codeword_reg5[256*9+2], codeword_reg4[256*9+2], codeword_reg3[256*9+2], codeword_reg2[256*9+2], codeword_reg1[256*9+2], codeword_reg16[256*8+2], codeword_reg15[256*8+2], codeword_reg14[256*8+2], codeword_reg13[256*8+2], codeword_reg12[256*8+2], codeword_reg11[256*8+2], codeword_reg10[256*8+2], codeword_reg9[256*8+2], codeword_reg8[256*8+2], codeword_reg7[256*8+2], codeword_reg6[256*8+2], codeword_reg5[256*8+2], codeword_reg4[256*8+2], codeword_reg3[256*8+2], codeword_reg2[256*8+2], codeword_reg1[256*8+2], codeword_reg16[256*7+2], codeword_reg15[256*7+2], codeword_reg14[256*7+2], codeword_reg13[256*7+2], codeword_reg12[256*7+2], codeword_reg11[256*7+2], codeword_reg10[256*7+2], codeword_reg9[256*7+2], codeword_reg8[256*7+2], codeword_reg7[256*7+2], codeword_reg6[256*7+2], codeword_reg5[256*7+2], codeword_reg4[256*7+2], codeword_reg3[256*7+2], codeword_reg2[256*7+2], codeword_reg1[256*7+2], codeword_reg16[256*6+2], codeword_reg15[256*6+2], codeword_reg14[256*6+2], codeword_reg13[256*6+2], codeword_reg12[256*6+2], codeword_reg11[256*6+2], codeword_reg10[256*6+2], codeword_reg9[256*6+2], codeword_reg8[256*6+2], codeword_reg7[256*6+2], codeword_reg6[256*6+2], codeword_reg5[256*6+2], codeword_reg4[256*6+2], codeword_reg3[256*6+2], codeword_reg2[256*6+2], codeword_reg1[256*6+2], codeword_reg16[256*5+2], codeword_reg15[256*5+2], codeword_reg14[256*5+2], codeword_reg13[256*5+2], codeword_reg12[256*5+2], codeword_reg11[256*5+2], codeword_reg10[256*5+2], codeword_reg9[256*5+2], codeword_reg8[256*5+2], codeword_reg7[256*5+2], codeword_reg6[256*5+2], codeword_reg5[256*5+2], codeword_reg4[256*5+2], codeword_reg3[256*5+2], codeword_reg2[256*5+2], codeword_reg1[256*5+2], codeword_reg16[256*4+2], codeword_reg15[256*4+2], codeword_reg14[256*4+2], codeword_reg13[256*4+2], codeword_reg12[256*4+2], codeword_reg11[256*4+2], codeword_reg10[256*4+2], codeword_reg9[256*4+2], codeword_reg8[256*4+2], codeword_reg7[256*4+2], codeword_reg6[256*4+2], codeword_reg5[256*4+2], codeword_reg4[256*4+2], codeword_reg3[256*4+2], codeword_reg2[256*4+2], codeword_reg1[256*4+2], codeword_reg16[256*3+2], codeword_reg15[256*3+2], codeword_reg14[256*3+2], codeword_reg13[256*3+2], codeword_reg12[256*3+2], codeword_reg11[256*3+2], codeword_reg10[256*3+2], codeword_reg9[256*3+2], codeword_reg8[256*3+2], codeword_reg7[256*3+2], codeword_reg6[256*3+2], codeword_reg5[256*3+2], codeword_reg4[256*3+2], codeword_reg3[256*3+2], codeword_reg2[256*3+2], codeword_reg1[256*3+2], codeword_reg16[256*2+2], codeword_reg15[256*2+2], codeword_reg14[256*2+2], codeword_reg13[256*2+2], codeword_reg12[256*2+2], codeword_reg11[256*2+2], codeword_reg10[256*2+2], codeword_reg9[256*2+2], codeword_reg8[256*2+2], codeword_reg7[256*2+2], codeword_reg6[256*2+2], codeword_reg5[256*2+2], codeword_reg4[256*2+2], codeword_reg3[256*2+2], codeword_reg2[256*2+2], codeword_reg1[256*2+2], codeword_reg16[256*1+2], codeword_reg15[256*1+2], codeword_reg14[256*1+2], codeword_reg13[256*1+2], codeword_reg12[256*1+2], codeword_reg11[256*1+2], codeword_reg10[256*1+2], codeword_reg9[256*1+2], codeword_reg8[256*1+2], codeword_reg7[256*1+2], codeword_reg6[256*1+2], codeword_reg5[256*1+2], codeword_reg4[256*1+2], codeword_reg3[256*1+2], codeword_reg2[256*1+2], codeword_reg1[256*1+2], codeword_reg16[256*0+2], codeword_reg15[256*0+2], codeword_reg14[256*0+2], codeword_reg13[256*0+2], codeword_reg12[256*0+2], codeword_reg11[256*0+2], codeword_reg10[256*0+2], codeword_reg9[256*0+2], codeword_reg8[256*0+2], codeword_reg7[256*0+2], codeword_reg6[256*0+2], codeword_reg5[256*0+2], codeword_reg4[256*0+2], codeword_reg3[256*0+2], codeword_reg2[256*0+2], codeword_reg1[256*0+2]};
                                in_bits4 <= {codeword16[3], codeword15[3], codeword14[3], codeword13[3], codeword12[3], codeword11[3], codeword10[3], codeword9[3], codeword8[3], codeword7[3], codeword6[3], codeword5[3], codeword4[3], codeword3[3], codeword2[3], codeword1[3], codeword_reg16[256*13+3], codeword_reg15[256*13+3], codeword_reg14[256*13+3], codeword_reg13[256*13+3], codeword_reg12[256*13+3], codeword_reg11[256*13+3], codeword_reg10[256*13+3], codeword_reg9[256*13+3], codeword_reg8[256*13+3], codeword_reg7[256*13+3], codeword_reg6[256*13+3], codeword_reg5[256*13+3], codeword_reg4[256*13+3], codeword_reg3[256*13+3], codeword_reg2[256*13+3], codeword_reg1[256*13+3], codeword_reg16[256*12+3], codeword_reg15[256*12+3], codeword_reg14[256*12+3], codeword_reg13[256*12+3], codeword_reg12[256*12+3], codeword_reg11[256*12+3], codeword_reg10[256*12+3], codeword_reg9[256*12+3], codeword_reg8[256*12+3], codeword_reg7[256*12+3], codeword_reg6[256*12+3], codeword_reg5[256*12+3], codeword_reg4[256*12+3], codeword_reg3[256*12+3], codeword_reg2[256*12+3], codeword_reg1[256*12+3], codeword_reg16[256*11+3], codeword_reg15[256*11+3], codeword_reg14[256*11+3], codeword_reg13[256*11+3], codeword_reg12[256*11+3], codeword_reg11[256*11+3], codeword_reg10[256*11+3], codeword_reg9[256*11+3], codeword_reg8[256*11+3], codeword_reg7[256*11+3], codeword_reg6[256*11+3], codeword_reg5[256*11+3], codeword_reg4[256*11+3], codeword_reg3[256*11+3], codeword_reg2[256*11+3], codeword_reg1[256*11+3], codeword_reg16[256*10+3], codeword_reg15[256*10+3], codeword_reg14[256*10+3], codeword_reg13[256*10+3], codeword_reg12[256*10+3], codeword_reg11[256*10+3], codeword_reg10[256*10+3], codeword_reg9[256*10+3], codeword_reg8[256*10+3], codeword_reg7[256*10+3], codeword_reg6[256*10+3], codeword_reg5[256*10+3], codeword_reg4[256*10+3], codeword_reg3[256*10+3], codeword_reg2[256*10+3], codeword_reg1[256*10+3], codeword_reg16[256*9+3], codeword_reg15[256*9+3], codeword_reg14[256*9+3], codeword_reg13[256*9+3], codeword_reg12[256*9+3], codeword_reg11[256*9+3], codeword_reg10[256*9+3], codeword_reg9[256*9+3], codeword_reg8[256*9+3], codeword_reg7[256*9+3], codeword_reg6[256*9+3], codeword_reg5[256*9+3], codeword_reg4[256*9+3], codeword_reg3[256*9+3], codeword_reg2[256*9+3], codeword_reg1[256*9+3], codeword_reg16[256*8+3], codeword_reg15[256*8+3], codeword_reg14[256*8+3], codeword_reg13[256*8+3], codeword_reg12[256*8+3], codeword_reg11[256*8+3], codeword_reg10[256*8+3], codeword_reg9[256*8+3], codeword_reg8[256*8+3], codeword_reg7[256*8+3], codeword_reg6[256*8+3], codeword_reg5[256*8+3], codeword_reg4[256*8+3], codeword_reg3[256*8+3], codeword_reg2[256*8+3], codeword_reg1[256*8+3], codeword_reg16[256*7+3], codeword_reg15[256*7+3], codeword_reg14[256*7+3], codeword_reg13[256*7+3], codeword_reg12[256*7+3], codeword_reg11[256*7+3], codeword_reg10[256*7+3], codeword_reg9[256*7+3], codeword_reg8[256*7+3], codeword_reg7[256*7+3], codeword_reg6[256*7+3], codeword_reg5[256*7+3], codeword_reg4[256*7+3], codeword_reg3[256*7+3], codeword_reg2[256*7+3], codeword_reg1[256*7+3], codeword_reg16[256*6+3], codeword_reg15[256*6+3], codeword_reg14[256*6+3], codeword_reg13[256*6+3], codeword_reg12[256*6+3], codeword_reg11[256*6+3], codeword_reg10[256*6+3], codeword_reg9[256*6+3], codeword_reg8[256*6+3], codeword_reg7[256*6+3], codeword_reg6[256*6+3], codeword_reg5[256*6+3], codeword_reg4[256*6+3], codeword_reg3[256*6+3], codeword_reg2[256*6+3], codeword_reg1[256*6+3], codeword_reg16[256*5+3], codeword_reg15[256*5+3], codeword_reg14[256*5+3], codeword_reg13[256*5+3], codeword_reg12[256*5+3], codeword_reg11[256*5+3], codeword_reg10[256*5+3], codeword_reg9[256*5+3], codeword_reg8[256*5+3], codeword_reg7[256*5+3], codeword_reg6[256*5+3], codeword_reg5[256*5+3], codeword_reg4[256*5+3], codeword_reg3[256*5+3], codeword_reg2[256*5+3], codeword_reg1[256*5+3], codeword_reg16[256*4+3], codeword_reg15[256*4+3], codeword_reg14[256*4+3], codeword_reg13[256*4+3], codeword_reg12[256*4+3], codeword_reg11[256*4+3], codeword_reg10[256*4+3], codeword_reg9[256*4+3], codeword_reg8[256*4+3], codeword_reg7[256*4+3], codeword_reg6[256*4+3], codeword_reg5[256*4+3], codeword_reg4[256*4+3], codeword_reg3[256*4+3], codeword_reg2[256*4+3], codeword_reg1[256*4+3], codeword_reg16[256*3+3], codeword_reg15[256*3+3], codeword_reg14[256*3+3], codeword_reg13[256*3+3], codeword_reg12[256*3+3], codeword_reg11[256*3+3], codeword_reg10[256*3+3], codeword_reg9[256*3+3], codeword_reg8[256*3+3], codeword_reg7[256*3+3], codeword_reg6[256*3+3], codeword_reg5[256*3+3], codeword_reg4[256*3+3], codeword_reg3[256*3+3], codeword_reg2[256*3+3], codeword_reg1[256*3+3], codeword_reg16[256*2+3], codeword_reg15[256*2+3], codeword_reg14[256*2+3], codeword_reg13[256*2+3], codeword_reg12[256*2+3], codeword_reg11[256*2+3], codeword_reg10[256*2+3], codeword_reg9[256*2+3], codeword_reg8[256*2+3], codeword_reg7[256*2+3], codeword_reg6[256*2+3], codeword_reg5[256*2+3], codeword_reg4[256*2+3], codeword_reg3[256*2+3], codeword_reg2[256*2+3], codeword_reg1[256*2+3], codeword_reg16[256*1+3], codeword_reg15[256*1+3], codeword_reg14[256*1+3], codeword_reg13[256*1+3], codeword_reg12[256*1+3], codeword_reg11[256*1+3], codeword_reg10[256*1+3], codeword_reg9[256*1+3], codeword_reg8[256*1+3], codeword_reg7[256*1+3], codeword_reg6[256*1+3], codeword_reg5[256*1+3], codeword_reg4[256*1+3], codeword_reg3[256*1+3], codeword_reg2[256*1+3], codeword_reg1[256*1+3], codeword_reg16[256*0+3], codeword_reg15[256*0+3], codeword_reg14[256*0+3], codeword_reg13[256*0+3], codeword_reg12[256*0+3], codeword_reg11[256*0+3], codeword_reg10[256*0+3], codeword_reg9[256*0+3], codeword_reg8[256*0+3], codeword_reg7[256*0+3], codeword_reg6[256*0+3], codeword_reg5[256*0+3], codeword_reg4[256*0+3], codeword_reg3[256*0+3], codeword_reg2[256*0+3], codeword_reg1[256*0+3]};
                                in_bits5 <= {codeword16[4], codeword15[4], codeword14[4], codeword13[4], codeword12[4], codeword11[4], codeword10[4], codeword9[4], codeword8[4], codeword7[4], codeword6[4], codeword5[4], codeword4[4], codeword3[4], codeword2[4], codeword1[4], codeword_reg16[256*13+4], codeword_reg15[256*13+4], codeword_reg14[256*13+4], codeword_reg13[256*13+4], codeword_reg12[256*13+4], codeword_reg11[256*13+4], codeword_reg10[256*13+4], codeword_reg9[256*13+4], codeword_reg8[256*13+4], codeword_reg7[256*13+4], codeword_reg6[256*13+4], codeword_reg5[256*13+4], codeword_reg4[256*13+4], codeword_reg3[256*13+4], codeword_reg2[256*13+4], codeword_reg1[256*13+4], codeword_reg16[256*12+4], codeword_reg15[256*12+4], codeword_reg14[256*12+4], codeword_reg13[256*12+4], codeword_reg12[256*12+4], codeword_reg11[256*12+4], codeword_reg10[256*12+4], codeword_reg9[256*12+4], codeword_reg8[256*12+4], codeword_reg7[256*12+4], codeword_reg6[256*12+4], codeword_reg5[256*12+4], codeword_reg4[256*12+4], codeword_reg3[256*12+4], codeword_reg2[256*12+4], codeword_reg1[256*12+4], codeword_reg16[256*11+4], codeword_reg15[256*11+4], codeword_reg14[256*11+4], codeword_reg13[256*11+4], codeword_reg12[256*11+4], codeword_reg11[256*11+4], codeword_reg10[256*11+4], codeword_reg9[256*11+4], codeword_reg8[256*11+4], codeword_reg7[256*11+4], codeword_reg6[256*11+4], codeword_reg5[256*11+4], codeword_reg4[256*11+4], codeword_reg3[256*11+4], codeword_reg2[256*11+4], codeword_reg1[256*11+4], codeword_reg16[256*10+4], codeword_reg15[256*10+4], codeword_reg14[256*10+4], codeword_reg13[256*10+4], codeword_reg12[256*10+4], codeword_reg11[256*10+4], codeword_reg10[256*10+4], codeword_reg9[256*10+4], codeword_reg8[256*10+4], codeword_reg7[256*10+4], codeword_reg6[256*10+4], codeword_reg5[256*10+4], codeword_reg4[256*10+4], codeword_reg3[256*10+4], codeword_reg2[256*10+4], codeword_reg1[256*10+4], codeword_reg16[256*9+4], codeword_reg15[256*9+4], codeword_reg14[256*9+4], codeword_reg13[256*9+4], codeword_reg12[256*9+4], codeword_reg11[256*9+4], codeword_reg10[256*9+4], codeword_reg9[256*9+4], codeword_reg8[256*9+4], codeword_reg7[256*9+4], codeword_reg6[256*9+4], codeword_reg5[256*9+4], codeword_reg4[256*9+4], codeword_reg3[256*9+4], codeword_reg2[256*9+4], codeword_reg1[256*9+4], codeword_reg16[256*8+4], codeword_reg15[256*8+4], codeword_reg14[256*8+4], codeword_reg13[256*8+4], codeword_reg12[256*8+4], codeword_reg11[256*8+4], codeword_reg10[256*8+4], codeword_reg9[256*8+4], codeword_reg8[256*8+4], codeword_reg7[256*8+4], codeword_reg6[256*8+4], codeword_reg5[256*8+4], codeword_reg4[256*8+4], codeword_reg3[256*8+4], codeword_reg2[256*8+4], codeword_reg1[256*8+4], codeword_reg16[256*7+4], codeword_reg15[256*7+4], codeword_reg14[256*7+4], codeword_reg13[256*7+4], codeword_reg12[256*7+4], codeword_reg11[256*7+4], codeword_reg10[256*7+4], codeword_reg9[256*7+4], codeword_reg8[256*7+4], codeword_reg7[256*7+4], codeword_reg6[256*7+4], codeword_reg5[256*7+4], codeword_reg4[256*7+4], codeword_reg3[256*7+4], codeword_reg2[256*7+4], codeword_reg1[256*7+4], codeword_reg16[256*6+4], codeword_reg15[256*6+4], codeword_reg14[256*6+4], codeword_reg13[256*6+4], codeword_reg12[256*6+4], codeword_reg11[256*6+4], codeword_reg10[256*6+4], codeword_reg9[256*6+4], codeword_reg8[256*6+4], codeword_reg7[256*6+4], codeword_reg6[256*6+4], codeword_reg5[256*6+4], codeword_reg4[256*6+4], codeword_reg3[256*6+4], codeword_reg2[256*6+4], codeword_reg1[256*6+4], codeword_reg16[256*5+4], codeword_reg15[256*5+4], codeword_reg14[256*5+4], codeword_reg13[256*5+4], codeword_reg12[256*5+4], codeword_reg11[256*5+4], codeword_reg10[256*5+4], codeword_reg9[256*5+4], codeword_reg8[256*5+4], codeword_reg7[256*5+4], codeword_reg6[256*5+4], codeword_reg5[256*5+4], codeword_reg4[256*5+4], codeword_reg3[256*5+4], codeword_reg2[256*5+4], codeword_reg1[256*5+4], codeword_reg16[256*4+4], codeword_reg15[256*4+4], codeword_reg14[256*4+4], codeword_reg13[256*4+4], codeword_reg12[256*4+4], codeword_reg11[256*4+4], codeword_reg10[256*4+4], codeword_reg9[256*4+4], codeword_reg8[256*4+4], codeword_reg7[256*4+4], codeword_reg6[256*4+4], codeword_reg5[256*4+4], codeword_reg4[256*4+4], codeword_reg3[256*4+4], codeword_reg2[256*4+4], codeword_reg1[256*4+4], codeword_reg16[256*3+4], codeword_reg15[256*3+4], codeword_reg14[256*3+4], codeword_reg13[256*3+4], codeword_reg12[256*3+4], codeword_reg11[256*3+4], codeword_reg10[256*3+4], codeword_reg9[256*3+4], codeword_reg8[256*3+4], codeword_reg7[256*3+4], codeword_reg6[256*3+4], codeword_reg5[256*3+4], codeword_reg4[256*3+4], codeword_reg3[256*3+4], codeword_reg2[256*3+4], codeword_reg1[256*3+4], codeword_reg16[256*2+4], codeword_reg15[256*2+4], codeword_reg14[256*2+4], codeword_reg13[256*2+4], codeword_reg12[256*2+4], codeword_reg11[256*2+4], codeword_reg10[256*2+4], codeword_reg9[256*2+4], codeword_reg8[256*2+4], codeword_reg7[256*2+4], codeword_reg6[256*2+4], codeword_reg5[256*2+4], codeword_reg4[256*2+4], codeword_reg3[256*2+4], codeword_reg2[256*2+4], codeword_reg1[256*2+4], codeword_reg16[256*1+4], codeword_reg15[256*1+4], codeword_reg14[256*1+4], codeword_reg13[256*1+4], codeword_reg12[256*1+4], codeword_reg11[256*1+4], codeword_reg10[256*1+4], codeword_reg9[256*1+4], codeword_reg8[256*1+4], codeword_reg7[256*1+4], codeword_reg6[256*1+4], codeword_reg5[256*1+4], codeword_reg4[256*1+4], codeword_reg3[256*1+4], codeword_reg2[256*1+4], codeword_reg1[256*1+4], codeword_reg16[256*0+4], codeword_reg15[256*0+4], codeword_reg14[256*0+4], codeword_reg13[256*0+4], codeword_reg12[256*0+4], codeword_reg11[256*0+4], codeword_reg10[256*0+4], codeword_reg9[256*0+4], codeword_reg8[256*0+4], codeword_reg7[256*0+4], codeword_reg6[256*0+4], codeword_reg5[256*0+4], codeword_reg4[256*0+4], codeword_reg3[256*0+4], codeword_reg2[256*0+4], codeword_reg1[256*0+4]};
                                in_bits6 <= {codeword16[5], codeword15[5], codeword14[5], codeword13[5], codeword12[5], codeword11[5], codeword10[5], codeword9[5], codeword8[5], codeword7[5], codeword6[5], codeword5[5], codeword4[5], codeword3[5], codeword2[5], codeword1[5], codeword_reg16[256*13+5], codeword_reg15[256*13+5], codeword_reg14[256*13+5], codeword_reg13[256*13+5], codeword_reg12[256*13+5], codeword_reg11[256*13+5], codeword_reg10[256*13+5], codeword_reg9[256*13+5], codeword_reg8[256*13+5], codeword_reg7[256*13+5], codeword_reg6[256*13+5], codeword_reg5[256*13+5], codeword_reg4[256*13+5], codeword_reg3[256*13+5], codeword_reg2[256*13+5], codeword_reg1[256*13+5], codeword_reg16[256*12+5], codeword_reg15[256*12+5], codeword_reg14[256*12+5], codeword_reg13[256*12+5], codeword_reg12[256*12+5], codeword_reg11[256*12+5], codeword_reg10[256*12+5], codeword_reg9[256*12+5], codeword_reg8[256*12+5], codeword_reg7[256*12+5], codeword_reg6[256*12+5], codeword_reg5[256*12+5], codeword_reg4[256*12+5], codeword_reg3[256*12+5], codeword_reg2[256*12+5], codeword_reg1[256*12+5], codeword_reg16[256*11+5], codeword_reg15[256*11+5], codeword_reg14[256*11+5], codeword_reg13[256*11+5], codeword_reg12[256*11+5], codeword_reg11[256*11+5], codeword_reg10[256*11+5], codeword_reg9[256*11+5], codeword_reg8[256*11+5], codeword_reg7[256*11+5], codeword_reg6[256*11+5], codeword_reg5[256*11+5], codeword_reg4[256*11+5], codeword_reg3[256*11+5], codeword_reg2[256*11+5], codeword_reg1[256*11+5], codeword_reg16[256*10+5], codeword_reg15[256*10+5], codeword_reg14[256*10+5], codeword_reg13[256*10+5], codeword_reg12[256*10+5], codeword_reg11[256*10+5], codeword_reg10[256*10+5], codeword_reg9[256*10+5], codeword_reg8[256*10+5], codeword_reg7[256*10+5], codeword_reg6[256*10+5], codeword_reg5[256*10+5], codeword_reg4[256*10+5], codeword_reg3[256*10+5], codeword_reg2[256*10+5], codeword_reg1[256*10+5], codeword_reg16[256*9+5], codeword_reg15[256*9+5], codeword_reg14[256*9+5], codeword_reg13[256*9+5], codeword_reg12[256*9+5], codeword_reg11[256*9+5], codeword_reg10[256*9+5], codeword_reg9[256*9+5], codeword_reg8[256*9+5], codeword_reg7[256*9+5], codeword_reg6[256*9+5], codeword_reg5[256*9+5], codeword_reg4[256*9+5], codeword_reg3[256*9+5], codeword_reg2[256*9+5], codeword_reg1[256*9+5], codeword_reg16[256*8+5], codeword_reg15[256*8+5], codeword_reg14[256*8+5], codeword_reg13[256*8+5], codeword_reg12[256*8+5], codeword_reg11[256*8+5], codeword_reg10[256*8+5], codeword_reg9[256*8+5], codeword_reg8[256*8+5], codeword_reg7[256*8+5], codeword_reg6[256*8+5], codeword_reg5[256*8+5], codeword_reg4[256*8+5], codeword_reg3[256*8+5], codeword_reg2[256*8+5], codeword_reg1[256*8+5], codeword_reg16[256*7+5], codeword_reg15[256*7+5], codeword_reg14[256*7+5], codeword_reg13[256*7+5], codeword_reg12[256*7+5], codeword_reg11[256*7+5], codeword_reg10[256*7+5], codeword_reg9[256*7+5], codeword_reg8[256*7+5], codeword_reg7[256*7+5], codeword_reg6[256*7+5], codeword_reg5[256*7+5], codeword_reg4[256*7+5], codeword_reg3[256*7+5], codeword_reg2[256*7+5], codeword_reg1[256*7+5], codeword_reg16[256*6+5], codeword_reg15[256*6+5], codeword_reg14[256*6+5], codeword_reg13[256*6+5], codeword_reg12[256*6+5], codeword_reg11[256*6+5], codeword_reg10[256*6+5], codeword_reg9[256*6+5], codeword_reg8[256*6+5], codeword_reg7[256*6+5], codeword_reg6[256*6+5], codeword_reg5[256*6+5], codeword_reg4[256*6+5], codeword_reg3[256*6+5], codeword_reg2[256*6+5], codeword_reg1[256*6+5], codeword_reg16[256*5+5], codeword_reg15[256*5+5], codeword_reg14[256*5+5], codeword_reg13[256*5+5], codeword_reg12[256*5+5], codeword_reg11[256*5+5], codeword_reg10[256*5+5], codeword_reg9[256*5+5], codeword_reg8[256*5+5], codeword_reg7[256*5+5], codeword_reg6[256*5+5], codeword_reg5[256*5+5], codeword_reg4[256*5+5], codeword_reg3[256*5+5], codeword_reg2[256*5+5], codeword_reg1[256*5+5], codeword_reg16[256*4+5], codeword_reg15[256*4+5], codeword_reg14[256*4+5], codeword_reg13[256*4+5], codeword_reg12[256*4+5], codeword_reg11[256*4+5], codeword_reg10[256*4+5], codeword_reg9[256*4+5], codeword_reg8[256*4+5], codeword_reg7[256*4+5], codeword_reg6[256*4+5], codeword_reg5[256*4+5], codeword_reg4[256*4+5], codeword_reg3[256*4+5], codeword_reg2[256*4+5], codeword_reg1[256*4+5], codeword_reg16[256*3+5], codeword_reg15[256*3+5], codeword_reg14[256*3+5], codeword_reg13[256*3+5], codeword_reg12[256*3+5], codeword_reg11[256*3+5], codeword_reg10[256*3+5], codeword_reg9[256*3+5], codeword_reg8[256*3+5], codeword_reg7[256*3+5], codeword_reg6[256*3+5], codeword_reg5[256*3+5], codeword_reg4[256*3+5], codeword_reg3[256*3+5], codeword_reg2[256*3+5], codeword_reg1[256*3+5], codeword_reg16[256*2+5], codeword_reg15[256*2+5], codeword_reg14[256*2+5], codeword_reg13[256*2+5], codeword_reg12[256*2+5], codeword_reg11[256*2+5], codeword_reg10[256*2+5], codeword_reg9[256*2+5], codeword_reg8[256*2+5], codeword_reg7[256*2+5], codeword_reg6[256*2+5], codeword_reg5[256*2+5], codeword_reg4[256*2+5], codeword_reg3[256*2+5], codeword_reg2[256*2+5], codeword_reg1[256*2+5], codeword_reg16[256*1+5], codeword_reg15[256*1+5], codeword_reg14[256*1+5], codeword_reg13[256*1+5], codeword_reg12[256*1+5], codeword_reg11[256*1+5], codeword_reg10[256*1+5], codeword_reg9[256*1+5], codeword_reg8[256*1+5], codeword_reg7[256*1+5], codeword_reg6[256*1+5], codeword_reg5[256*1+5], codeword_reg4[256*1+5], codeword_reg3[256*1+5], codeword_reg2[256*1+5], codeword_reg1[256*1+5], codeword_reg16[256*0+5], codeword_reg15[256*0+5], codeword_reg14[256*0+5], codeword_reg13[256*0+5], codeword_reg12[256*0+5], codeword_reg11[256*0+5], codeword_reg10[256*0+5], codeword_reg9[256*0+5], codeword_reg8[256*0+5], codeword_reg7[256*0+5], codeword_reg6[256*0+5], codeword_reg5[256*0+5], codeword_reg4[256*0+5], codeword_reg3[256*0+5], codeword_reg2[256*0+5], codeword_reg1[256*0+5]};
                                in_bits7 <= {codeword16[6], codeword15[6], codeword14[6], codeword13[6], codeword12[6], codeword11[6], codeword10[6], codeword9[6], codeword8[6], codeword7[6], codeword6[6], codeword5[6], codeword4[6], codeword3[6], codeword2[6], codeword1[6], codeword_reg16[256*13+6], codeword_reg15[256*13+6], codeword_reg14[256*13+6], codeword_reg13[256*13+6], codeword_reg12[256*13+6], codeword_reg11[256*13+6], codeword_reg10[256*13+6], codeword_reg9[256*13+6], codeword_reg8[256*13+6], codeword_reg7[256*13+6], codeword_reg6[256*13+6], codeword_reg5[256*13+6], codeword_reg4[256*13+6], codeword_reg3[256*13+6], codeword_reg2[256*13+6], codeword_reg1[256*13+6], codeword_reg16[256*12+6], codeword_reg15[256*12+6], codeword_reg14[256*12+6], codeword_reg13[256*12+6], codeword_reg12[256*12+6], codeword_reg11[256*12+6], codeword_reg10[256*12+6], codeword_reg9[256*12+6], codeword_reg8[256*12+6], codeword_reg7[256*12+6], codeword_reg6[256*12+6], codeword_reg5[256*12+6], codeword_reg4[256*12+6], codeword_reg3[256*12+6], codeword_reg2[256*12+6], codeword_reg1[256*12+6], codeword_reg16[256*11+6], codeword_reg15[256*11+6], codeword_reg14[256*11+6], codeword_reg13[256*11+6], codeword_reg12[256*11+6], codeword_reg11[256*11+6], codeword_reg10[256*11+6], codeword_reg9[256*11+6], codeword_reg8[256*11+6], codeword_reg7[256*11+6], codeword_reg6[256*11+6], codeword_reg5[256*11+6], codeword_reg4[256*11+6], codeword_reg3[256*11+6], codeword_reg2[256*11+6], codeword_reg1[256*11+6], codeword_reg16[256*10+6], codeword_reg15[256*10+6], codeword_reg14[256*10+6], codeword_reg13[256*10+6], codeword_reg12[256*10+6], codeword_reg11[256*10+6], codeword_reg10[256*10+6], codeword_reg9[256*10+6], codeword_reg8[256*10+6], codeword_reg7[256*10+6], codeword_reg6[256*10+6], codeword_reg5[256*10+6], codeword_reg4[256*10+6], codeword_reg3[256*10+6], codeword_reg2[256*10+6], codeword_reg1[256*10+6], codeword_reg16[256*9+6], codeword_reg15[256*9+6], codeword_reg14[256*9+6], codeword_reg13[256*9+6], codeword_reg12[256*9+6], codeword_reg11[256*9+6], codeword_reg10[256*9+6], codeword_reg9[256*9+6], codeword_reg8[256*9+6], codeword_reg7[256*9+6], codeword_reg6[256*9+6], codeword_reg5[256*9+6], codeword_reg4[256*9+6], codeword_reg3[256*9+6], codeword_reg2[256*9+6], codeword_reg1[256*9+6], codeword_reg16[256*8+6], codeword_reg15[256*8+6], codeword_reg14[256*8+6], codeword_reg13[256*8+6], codeword_reg12[256*8+6], codeword_reg11[256*8+6], codeword_reg10[256*8+6], codeword_reg9[256*8+6], codeword_reg8[256*8+6], codeword_reg7[256*8+6], codeword_reg6[256*8+6], codeword_reg5[256*8+6], codeword_reg4[256*8+6], codeword_reg3[256*8+6], codeword_reg2[256*8+6], codeword_reg1[256*8+6], codeword_reg16[256*7+6], codeword_reg15[256*7+6], codeword_reg14[256*7+6], codeword_reg13[256*7+6], codeword_reg12[256*7+6], codeword_reg11[256*7+6], codeword_reg10[256*7+6], codeword_reg9[256*7+6], codeword_reg8[256*7+6], codeword_reg7[256*7+6], codeword_reg6[256*7+6], codeword_reg5[256*7+6], codeword_reg4[256*7+6], codeword_reg3[256*7+6], codeword_reg2[256*7+6], codeword_reg1[256*7+6], codeword_reg16[256*6+6], codeword_reg15[256*6+6], codeword_reg14[256*6+6], codeword_reg13[256*6+6], codeword_reg12[256*6+6], codeword_reg11[256*6+6], codeword_reg10[256*6+6], codeword_reg9[256*6+6], codeword_reg8[256*6+6], codeword_reg7[256*6+6], codeword_reg6[256*6+6], codeword_reg5[256*6+6], codeword_reg4[256*6+6], codeword_reg3[256*6+6], codeword_reg2[256*6+6], codeword_reg1[256*6+6], codeword_reg16[256*5+6], codeword_reg15[256*5+6], codeword_reg14[256*5+6], codeword_reg13[256*5+6], codeword_reg12[256*5+6], codeword_reg11[256*5+6], codeword_reg10[256*5+6], codeword_reg9[256*5+6], codeword_reg8[256*5+6], codeword_reg7[256*5+6], codeword_reg6[256*5+6], codeword_reg5[256*5+6], codeword_reg4[256*5+6], codeword_reg3[256*5+6], codeword_reg2[256*5+6], codeword_reg1[256*5+6], codeword_reg16[256*4+6], codeword_reg15[256*4+6], codeword_reg14[256*4+6], codeword_reg13[256*4+6], codeword_reg12[256*4+6], codeword_reg11[256*4+6], codeword_reg10[256*4+6], codeword_reg9[256*4+6], codeword_reg8[256*4+6], codeword_reg7[256*4+6], codeword_reg6[256*4+6], codeword_reg5[256*4+6], codeword_reg4[256*4+6], codeword_reg3[256*4+6], codeword_reg2[256*4+6], codeword_reg1[256*4+6], codeword_reg16[256*3+6], codeword_reg15[256*3+6], codeword_reg14[256*3+6], codeword_reg13[256*3+6], codeword_reg12[256*3+6], codeword_reg11[256*3+6], codeword_reg10[256*3+6], codeword_reg9[256*3+6], codeword_reg8[256*3+6], codeword_reg7[256*3+6], codeword_reg6[256*3+6], codeword_reg5[256*3+6], codeword_reg4[256*3+6], codeword_reg3[256*3+6], codeword_reg2[256*3+6], codeword_reg1[256*3+6], codeword_reg16[256*2+6], codeword_reg15[256*2+6], codeword_reg14[256*2+6], codeword_reg13[256*2+6], codeword_reg12[256*2+6], codeword_reg11[256*2+6], codeword_reg10[256*2+6], codeword_reg9[256*2+6], codeword_reg8[256*2+6], codeword_reg7[256*2+6], codeword_reg6[256*2+6], codeword_reg5[256*2+6], codeword_reg4[256*2+6], codeword_reg3[256*2+6], codeword_reg2[256*2+6], codeword_reg1[256*2+6], codeword_reg16[256*1+6], codeword_reg15[256*1+6], codeword_reg14[256*1+6], codeword_reg13[256*1+6], codeword_reg12[256*1+6], codeword_reg11[256*1+6], codeword_reg10[256*1+6], codeword_reg9[256*1+6], codeword_reg8[256*1+6], codeword_reg7[256*1+6], codeword_reg6[256*1+6], codeword_reg5[256*1+6], codeword_reg4[256*1+6], codeword_reg3[256*1+6], codeword_reg2[256*1+6], codeword_reg1[256*1+6], codeword_reg16[256*0+6], codeword_reg15[256*0+6], codeword_reg14[256*0+6], codeword_reg13[256*0+6], codeword_reg12[256*0+6], codeword_reg11[256*0+6], codeword_reg10[256*0+6], codeword_reg9[256*0+6], codeword_reg8[256*0+6], codeword_reg7[256*0+6], codeword_reg6[256*0+6], codeword_reg5[256*0+6], codeword_reg4[256*0+6], codeword_reg3[256*0+6], codeword_reg2[256*0+6], codeword_reg1[256*0+6]};
                                in_bits8 <= {codeword16[7], codeword15[7], codeword14[7], codeword13[7], codeword12[7], codeword11[7], codeword10[7], codeword9[7], codeword8[7], codeword7[7], codeword6[7], codeword5[7], codeword4[7], codeword3[7], codeword2[7], codeword1[7], codeword_reg16[256*13+7], codeword_reg15[256*13+7], codeword_reg14[256*13+7], codeword_reg13[256*13+7], codeword_reg12[256*13+7], codeword_reg11[256*13+7], codeword_reg10[256*13+7], codeword_reg9[256*13+7], codeword_reg8[256*13+7], codeword_reg7[256*13+7], codeword_reg6[256*13+7], codeword_reg5[256*13+7], codeword_reg4[256*13+7], codeword_reg3[256*13+7], codeword_reg2[256*13+7], codeword_reg1[256*13+7], codeword_reg16[256*12+7], codeword_reg15[256*12+7], codeword_reg14[256*12+7], codeword_reg13[256*12+7], codeword_reg12[256*12+7], codeword_reg11[256*12+7], codeword_reg10[256*12+7], codeword_reg9[256*12+7], codeword_reg8[256*12+7], codeword_reg7[256*12+7], codeword_reg6[256*12+7], codeword_reg5[256*12+7], codeword_reg4[256*12+7], codeword_reg3[256*12+7], codeword_reg2[256*12+7], codeword_reg1[256*12+7], codeword_reg16[256*11+7], codeword_reg15[256*11+7], codeword_reg14[256*11+7], codeword_reg13[256*11+7], codeword_reg12[256*11+7], codeword_reg11[256*11+7], codeword_reg10[256*11+7], codeword_reg9[256*11+7], codeword_reg8[256*11+7], codeword_reg7[256*11+7], codeword_reg6[256*11+7], codeword_reg5[256*11+7], codeword_reg4[256*11+7], codeword_reg3[256*11+7], codeword_reg2[256*11+7], codeword_reg1[256*11+7], codeword_reg16[256*10+7], codeword_reg15[256*10+7], codeword_reg14[256*10+7], codeword_reg13[256*10+7], codeword_reg12[256*10+7], codeword_reg11[256*10+7], codeword_reg10[256*10+7], codeword_reg9[256*10+7], codeword_reg8[256*10+7], codeword_reg7[256*10+7], codeword_reg6[256*10+7], codeword_reg5[256*10+7], codeword_reg4[256*10+7], codeword_reg3[256*10+7], codeword_reg2[256*10+7], codeword_reg1[256*10+7], codeword_reg16[256*9+7], codeword_reg15[256*9+7], codeword_reg14[256*9+7], codeword_reg13[256*9+7], codeword_reg12[256*9+7], codeword_reg11[256*9+7], codeword_reg10[256*9+7], codeword_reg9[256*9+7], codeword_reg8[256*9+7], codeword_reg7[256*9+7], codeword_reg6[256*9+7], codeword_reg5[256*9+7], codeword_reg4[256*9+7], codeword_reg3[256*9+7], codeword_reg2[256*9+7], codeword_reg1[256*9+7], codeword_reg16[256*8+7], codeword_reg15[256*8+7], codeword_reg14[256*8+7], codeword_reg13[256*8+7], codeword_reg12[256*8+7], codeword_reg11[256*8+7], codeword_reg10[256*8+7], codeword_reg9[256*8+7], codeword_reg8[256*8+7], codeword_reg7[256*8+7], codeword_reg6[256*8+7], codeword_reg5[256*8+7], codeword_reg4[256*8+7], codeword_reg3[256*8+7], codeword_reg2[256*8+7], codeword_reg1[256*8+7], codeword_reg16[256*7+7], codeword_reg15[256*7+7], codeword_reg14[256*7+7], codeword_reg13[256*7+7], codeword_reg12[256*7+7], codeword_reg11[256*7+7], codeword_reg10[256*7+7], codeword_reg9[256*7+7], codeword_reg8[256*7+7], codeword_reg7[256*7+7], codeword_reg6[256*7+7], codeword_reg5[256*7+7], codeword_reg4[256*7+7], codeword_reg3[256*7+7], codeword_reg2[256*7+7], codeword_reg1[256*7+7], codeword_reg16[256*6+7], codeword_reg15[256*6+7], codeword_reg14[256*6+7], codeword_reg13[256*6+7], codeword_reg12[256*6+7], codeword_reg11[256*6+7], codeword_reg10[256*6+7], codeword_reg9[256*6+7], codeword_reg8[256*6+7], codeword_reg7[256*6+7], codeword_reg6[256*6+7], codeword_reg5[256*6+7], codeword_reg4[256*6+7], codeword_reg3[256*6+7], codeword_reg2[256*6+7], codeword_reg1[256*6+7], codeword_reg16[256*5+7], codeword_reg15[256*5+7], codeword_reg14[256*5+7], codeword_reg13[256*5+7], codeword_reg12[256*5+7], codeword_reg11[256*5+7], codeword_reg10[256*5+7], codeword_reg9[256*5+7], codeword_reg8[256*5+7], codeword_reg7[256*5+7], codeword_reg6[256*5+7], codeword_reg5[256*5+7], codeword_reg4[256*5+7], codeword_reg3[256*5+7], codeword_reg2[256*5+7], codeword_reg1[256*5+7], codeword_reg16[256*4+7], codeword_reg15[256*4+7], codeword_reg14[256*4+7], codeword_reg13[256*4+7], codeword_reg12[256*4+7], codeword_reg11[256*4+7], codeword_reg10[256*4+7], codeword_reg9[256*4+7], codeword_reg8[256*4+7], codeword_reg7[256*4+7], codeword_reg6[256*4+7], codeword_reg5[256*4+7], codeword_reg4[256*4+7], codeword_reg3[256*4+7], codeword_reg2[256*4+7], codeword_reg1[256*4+7], codeword_reg16[256*3+7], codeword_reg15[256*3+7], codeword_reg14[256*3+7], codeword_reg13[256*3+7], codeword_reg12[256*3+7], codeword_reg11[256*3+7], codeword_reg10[256*3+7], codeword_reg9[256*3+7], codeword_reg8[256*3+7], codeword_reg7[256*3+7], codeword_reg6[256*3+7], codeword_reg5[256*3+7], codeword_reg4[256*3+7], codeword_reg3[256*3+7], codeword_reg2[256*3+7], codeword_reg1[256*3+7], codeword_reg16[256*2+7], codeword_reg15[256*2+7], codeword_reg14[256*2+7], codeword_reg13[256*2+7], codeword_reg12[256*2+7], codeword_reg11[256*2+7], codeword_reg10[256*2+7], codeword_reg9[256*2+7], codeword_reg8[256*2+7], codeword_reg7[256*2+7], codeword_reg6[256*2+7], codeword_reg5[256*2+7], codeword_reg4[256*2+7], codeword_reg3[256*2+7], codeword_reg2[256*2+7], codeword_reg1[256*2+7], codeword_reg16[256*1+7], codeword_reg15[256*1+7], codeword_reg14[256*1+7], codeword_reg13[256*1+7], codeword_reg12[256*1+7], codeword_reg11[256*1+7], codeword_reg10[256*1+7], codeword_reg9[256*1+7], codeword_reg8[256*1+7], codeword_reg7[256*1+7], codeword_reg6[256*1+7], codeword_reg5[256*1+7], codeword_reg4[256*1+7], codeword_reg3[256*1+7], codeword_reg2[256*1+7], codeword_reg1[256*1+7], codeword_reg16[256*0+7], codeword_reg15[256*0+7], codeword_reg14[256*0+7], codeword_reg13[256*0+7], codeword_reg12[256*0+7], codeword_reg11[256*0+7], codeword_reg10[256*0+7], codeword_reg9[256*0+7], codeword_reg8[256*0+7], codeword_reg7[256*0+7], codeword_reg6[256*0+7], codeword_reg5[256*0+7], codeword_reg4[256*0+7], codeword_reg3[256*0+7], codeword_reg2[256*0+7], codeword_reg1[256*0+7]};
                                in_bits9 <= {codeword16[8], codeword15[8], codeword14[8], codeword13[8], codeword12[8], codeword11[8], codeword10[8], codeword9[8], codeword8[8], codeword7[8], codeword6[8], codeword5[8], codeword4[8], codeword3[8], codeword2[8], codeword1[8], codeword_reg16[256*13+8], codeword_reg15[256*13+8], codeword_reg14[256*13+8], codeword_reg13[256*13+8], codeword_reg12[256*13+8], codeword_reg11[256*13+8], codeword_reg10[256*13+8], codeword_reg9[256*13+8], codeword_reg8[256*13+8], codeword_reg7[256*13+8], codeword_reg6[256*13+8], codeword_reg5[256*13+8], codeword_reg4[256*13+8], codeword_reg3[256*13+8], codeword_reg2[256*13+8], codeword_reg1[256*13+8], codeword_reg16[256*12+8], codeword_reg15[256*12+8], codeword_reg14[256*12+8], codeword_reg13[256*12+8], codeword_reg12[256*12+8], codeword_reg11[256*12+8], codeword_reg10[256*12+8], codeword_reg9[256*12+8], codeword_reg8[256*12+8], codeword_reg7[256*12+8], codeword_reg6[256*12+8], codeword_reg5[256*12+8], codeword_reg4[256*12+8], codeword_reg3[256*12+8], codeword_reg2[256*12+8], codeword_reg1[256*12+8], codeword_reg16[256*11+8], codeword_reg15[256*11+8], codeword_reg14[256*11+8], codeword_reg13[256*11+8], codeword_reg12[256*11+8], codeword_reg11[256*11+8], codeword_reg10[256*11+8], codeword_reg9[256*11+8], codeword_reg8[256*11+8], codeword_reg7[256*11+8], codeword_reg6[256*11+8], codeword_reg5[256*11+8], codeword_reg4[256*11+8], codeword_reg3[256*11+8], codeword_reg2[256*11+8], codeword_reg1[256*11+8], codeword_reg16[256*10+8], codeword_reg15[256*10+8], codeword_reg14[256*10+8], codeword_reg13[256*10+8], codeword_reg12[256*10+8], codeword_reg11[256*10+8], codeword_reg10[256*10+8], codeword_reg9[256*10+8], codeword_reg8[256*10+8], codeword_reg7[256*10+8], codeword_reg6[256*10+8], codeword_reg5[256*10+8], codeword_reg4[256*10+8], codeword_reg3[256*10+8], codeword_reg2[256*10+8], codeword_reg1[256*10+8], codeword_reg16[256*9+8], codeword_reg15[256*9+8], codeword_reg14[256*9+8], codeword_reg13[256*9+8], codeword_reg12[256*9+8], codeword_reg11[256*9+8], codeword_reg10[256*9+8], codeword_reg9[256*9+8], codeword_reg8[256*9+8], codeword_reg7[256*9+8], codeword_reg6[256*9+8], codeword_reg5[256*9+8], codeword_reg4[256*9+8], codeword_reg3[256*9+8], codeword_reg2[256*9+8], codeword_reg1[256*9+8], codeword_reg16[256*8+8], codeword_reg15[256*8+8], codeword_reg14[256*8+8], codeword_reg13[256*8+8], codeword_reg12[256*8+8], codeword_reg11[256*8+8], codeword_reg10[256*8+8], codeword_reg9[256*8+8], codeword_reg8[256*8+8], codeword_reg7[256*8+8], codeword_reg6[256*8+8], codeword_reg5[256*8+8], codeword_reg4[256*8+8], codeword_reg3[256*8+8], codeword_reg2[256*8+8], codeword_reg1[256*8+8], codeword_reg16[256*7+8], codeword_reg15[256*7+8], codeword_reg14[256*7+8], codeword_reg13[256*7+8], codeword_reg12[256*7+8], codeword_reg11[256*7+8], codeword_reg10[256*7+8], codeword_reg9[256*7+8], codeword_reg8[256*7+8], codeword_reg7[256*7+8], codeword_reg6[256*7+8], codeword_reg5[256*7+8], codeword_reg4[256*7+8], codeword_reg3[256*7+8], codeword_reg2[256*7+8], codeword_reg1[256*7+8], codeword_reg16[256*6+8], codeword_reg15[256*6+8], codeword_reg14[256*6+8], codeword_reg13[256*6+8], codeword_reg12[256*6+8], codeword_reg11[256*6+8], codeword_reg10[256*6+8], codeword_reg9[256*6+8], codeword_reg8[256*6+8], codeword_reg7[256*6+8], codeword_reg6[256*6+8], codeword_reg5[256*6+8], codeword_reg4[256*6+8], codeword_reg3[256*6+8], codeword_reg2[256*6+8], codeword_reg1[256*6+8], codeword_reg16[256*5+8], codeword_reg15[256*5+8], codeword_reg14[256*5+8], codeword_reg13[256*5+8], codeword_reg12[256*5+8], codeword_reg11[256*5+8], codeword_reg10[256*5+8], codeword_reg9[256*5+8], codeword_reg8[256*5+8], codeword_reg7[256*5+8], codeword_reg6[256*5+8], codeword_reg5[256*5+8], codeword_reg4[256*5+8], codeword_reg3[256*5+8], codeword_reg2[256*5+8], codeword_reg1[256*5+8], codeword_reg16[256*4+8], codeword_reg15[256*4+8], codeword_reg14[256*4+8], codeword_reg13[256*4+8], codeword_reg12[256*4+8], codeword_reg11[256*4+8], codeword_reg10[256*4+8], codeword_reg9[256*4+8], codeword_reg8[256*4+8], codeword_reg7[256*4+8], codeword_reg6[256*4+8], codeword_reg5[256*4+8], codeword_reg4[256*4+8], codeword_reg3[256*4+8], codeword_reg2[256*4+8], codeword_reg1[256*4+8], codeword_reg16[256*3+8], codeword_reg15[256*3+8], codeword_reg14[256*3+8], codeword_reg13[256*3+8], codeword_reg12[256*3+8], codeword_reg11[256*3+8], codeword_reg10[256*3+8], codeword_reg9[256*3+8], codeword_reg8[256*3+8], codeword_reg7[256*3+8], codeword_reg6[256*3+8], codeword_reg5[256*3+8], codeword_reg4[256*3+8], codeword_reg3[256*3+8], codeword_reg2[256*3+8], codeword_reg1[256*3+8], codeword_reg16[256*2+8], codeword_reg15[256*2+8], codeword_reg14[256*2+8], codeword_reg13[256*2+8], codeword_reg12[256*2+8], codeword_reg11[256*2+8], codeword_reg10[256*2+8], codeword_reg9[256*2+8], codeword_reg8[256*2+8], codeword_reg7[256*2+8], codeword_reg6[256*2+8], codeword_reg5[256*2+8], codeword_reg4[256*2+8], codeword_reg3[256*2+8], codeword_reg2[256*2+8], codeword_reg1[256*2+8], codeword_reg16[256*1+8], codeword_reg15[256*1+8], codeword_reg14[256*1+8], codeword_reg13[256*1+8], codeword_reg12[256*1+8], codeword_reg11[256*1+8], codeword_reg10[256*1+8], codeword_reg9[256*1+8], codeword_reg8[256*1+8], codeword_reg7[256*1+8], codeword_reg6[256*1+8], codeword_reg5[256*1+8], codeword_reg4[256*1+8], codeword_reg3[256*1+8], codeword_reg2[256*1+8], codeword_reg1[256*1+8], codeword_reg16[256*0+8], codeword_reg15[256*0+8], codeword_reg14[256*0+8], codeword_reg13[256*0+8], codeword_reg12[256*0+8], codeword_reg11[256*0+8], codeword_reg10[256*0+8], codeword_reg9[256*0+8], codeword_reg8[256*0+8], codeword_reg7[256*0+8], codeword_reg6[256*0+8], codeword_reg5[256*0+8], codeword_reg4[256*0+8], codeword_reg3[256*0+8], codeword_reg2[256*0+8], codeword_reg1[256*0+8]};
                                in_bits10 <= {codeword16[9], codeword15[9], codeword14[9], codeword13[9], codeword12[9], codeword11[9], codeword10[9], codeword9[9], codeword8[9], codeword7[9], codeword6[9], codeword5[9], codeword4[9], codeword3[9], codeword2[9], codeword1[9], codeword_reg16[256*13+9], codeword_reg15[256*13+9], codeword_reg14[256*13+9], codeword_reg13[256*13+9], codeword_reg12[256*13+9], codeword_reg11[256*13+9], codeword_reg10[256*13+9], codeword_reg9[256*13+9], codeword_reg8[256*13+9], codeword_reg7[256*13+9], codeword_reg6[256*13+9], codeword_reg5[256*13+9], codeword_reg4[256*13+9], codeword_reg3[256*13+9], codeword_reg2[256*13+9], codeword_reg1[256*13+9], codeword_reg16[256*12+9], codeword_reg15[256*12+9], codeword_reg14[256*12+9], codeword_reg13[256*12+9], codeword_reg12[256*12+9], codeword_reg11[256*12+9], codeword_reg10[256*12+9], codeword_reg9[256*12+9], codeword_reg8[256*12+9], codeword_reg7[256*12+9], codeword_reg6[256*12+9], codeword_reg5[256*12+9], codeword_reg4[256*12+9], codeword_reg3[256*12+9], codeword_reg2[256*12+9], codeword_reg1[256*12+9], codeword_reg16[256*11+9], codeword_reg15[256*11+9], codeword_reg14[256*11+9], codeword_reg13[256*11+9], codeword_reg12[256*11+9], codeword_reg11[256*11+9], codeword_reg10[256*11+9], codeword_reg9[256*11+9], codeword_reg8[256*11+9], codeword_reg7[256*11+9], codeword_reg6[256*11+9], codeword_reg5[256*11+9], codeword_reg4[256*11+9], codeword_reg3[256*11+9], codeword_reg2[256*11+9], codeword_reg1[256*11+9], codeword_reg16[256*10+9], codeword_reg15[256*10+9], codeword_reg14[256*10+9], codeword_reg13[256*10+9], codeword_reg12[256*10+9], codeword_reg11[256*10+9], codeword_reg10[256*10+9], codeword_reg9[256*10+9], codeword_reg8[256*10+9], codeword_reg7[256*10+9], codeword_reg6[256*10+9], codeword_reg5[256*10+9], codeword_reg4[256*10+9], codeword_reg3[256*10+9], codeword_reg2[256*10+9], codeword_reg1[256*10+9], codeword_reg16[256*9+9], codeword_reg15[256*9+9], codeword_reg14[256*9+9], codeword_reg13[256*9+9], codeword_reg12[256*9+9], codeword_reg11[256*9+9], codeword_reg10[256*9+9], codeword_reg9[256*9+9], codeword_reg8[256*9+9], codeword_reg7[256*9+9], codeword_reg6[256*9+9], codeword_reg5[256*9+9], codeword_reg4[256*9+9], codeword_reg3[256*9+9], codeword_reg2[256*9+9], codeword_reg1[256*9+9], codeword_reg16[256*8+9], codeword_reg15[256*8+9], codeword_reg14[256*8+9], codeword_reg13[256*8+9], codeword_reg12[256*8+9], codeword_reg11[256*8+9], codeword_reg10[256*8+9], codeword_reg9[256*8+9], codeword_reg8[256*8+9], codeword_reg7[256*8+9], codeword_reg6[256*8+9], codeword_reg5[256*8+9], codeword_reg4[256*8+9], codeword_reg3[256*8+9], codeword_reg2[256*8+9], codeword_reg1[256*8+9], codeword_reg16[256*7+9], codeword_reg15[256*7+9], codeword_reg14[256*7+9], codeword_reg13[256*7+9], codeword_reg12[256*7+9], codeword_reg11[256*7+9], codeword_reg10[256*7+9], codeword_reg9[256*7+9], codeword_reg8[256*7+9], codeword_reg7[256*7+9], codeword_reg6[256*7+9], codeword_reg5[256*7+9], codeword_reg4[256*7+9], codeword_reg3[256*7+9], codeword_reg2[256*7+9], codeword_reg1[256*7+9], codeword_reg16[256*6+9], codeword_reg15[256*6+9], codeword_reg14[256*6+9], codeword_reg13[256*6+9], codeword_reg12[256*6+9], codeword_reg11[256*6+9], codeword_reg10[256*6+9], codeword_reg9[256*6+9], codeword_reg8[256*6+9], codeword_reg7[256*6+9], codeword_reg6[256*6+9], codeword_reg5[256*6+9], codeword_reg4[256*6+9], codeword_reg3[256*6+9], codeword_reg2[256*6+9], codeword_reg1[256*6+9], codeword_reg16[256*5+9], codeword_reg15[256*5+9], codeword_reg14[256*5+9], codeword_reg13[256*5+9], codeword_reg12[256*5+9], codeword_reg11[256*5+9], codeword_reg10[256*5+9], codeword_reg9[256*5+9], codeword_reg8[256*5+9], codeword_reg7[256*5+9], codeword_reg6[256*5+9], codeword_reg5[256*5+9], codeword_reg4[256*5+9], codeword_reg3[256*5+9], codeword_reg2[256*5+9], codeword_reg1[256*5+9], codeword_reg16[256*4+9], codeword_reg15[256*4+9], codeword_reg14[256*4+9], codeword_reg13[256*4+9], codeword_reg12[256*4+9], codeword_reg11[256*4+9], codeword_reg10[256*4+9], codeword_reg9[256*4+9], codeword_reg8[256*4+9], codeword_reg7[256*4+9], codeword_reg6[256*4+9], codeword_reg5[256*4+9], codeword_reg4[256*4+9], codeword_reg3[256*4+9], codeword_reg2[256*4+9], codeword_reg1[256*4+9], codeword_reg16[256*3+9], codeword_reg15[256*3+9], codeword_reg14[256*3+9], codeword_reg13[256*3+9], codeword_reg12[256*3+9], codeword_reg11[256*3+9], codeword_reg10[256*3+9], codeword_reg9[256*3+9], codeword_reg8[256*3+9], codeword_reg7[256*3+9], codeword_reg6[256*3+9], codeword_reg5[256*3+9], codeword_reg4[256*3+9], codeword_reg3[256*3+9], codeword_reg2[256*3+9], codeword_reg1[256*3+9], codeword_reg16[256*2+9], codeword_reg15[256*2+9], codeword_reg14[256*2+9], codeword_reg13[256*2+9], codeword_reg12[256*2+9], codeword_reg11[256*2+9], codeword_reg10[256*2+9], codeword_reg9[256*2+9], codeword_reg8[256*2+9], codeword_reg7[256*2+9], codeword_reg6[256*2+9], codeword_reg5[256*2+9], codeword_reg4[256*2+9], codeword_reg3[256*2+9], codeword_reg2[256*2+9], codeword_reg1[256*2+9], codeword_reg16[256*1+9], codeword_reg15[256*1+9], codeword_reg14[256*1+9], codeword_reg13[256*1+9], codeword_reg12[256*1+9], codeword_reg11[256*1+9], codeword_reg10[256*1+9], codeword_reg9[256*1+9], codeword_reg8[256*1+9], codeword_reg7[256*1+9], codeword_reg6[256*1+9], codeword_reg5[256*1+9], codeword_reg4[256*1+9], codeword_reg3[256*1+9], codeword_reg2[256*1+9], codeword_reg1[256*1+9], codeword_reg16[256*0+9], codeword_reg15[256*0+9], codeword_reg14[256*0+9], codeword_reg13[256*0+9], codeword_reg12[256*0+9], codeword_reg11[256*0+9], codeword_reg10[256*0+9], codeword_reg9[256*0+9], codeword_reg8[256*0+9], codeword_reg7[256*0+9], codeword_reg6[256*0+9], codeword_reg5[256*0+9], codeword_reg4[256*0+9], codeword_reg3[256*0+9], codeword_reg2[256*0+9], codeword_reg1[256*0+9]};
                                in_bits11 <= {codeword16[10], codeword15[10], codeword14[10], codeword13[10], codeword12[10], codeword11[10], codeword10[10], codeword9[10], codeword8[10], codeword7[10], codeword6[10], codeword5[10], codeword4[10], codeword3[10], codeword2[10], codeword1[10], codeword_reg16[256*13+10], codeword_reg15[256*13+10], codeword_reg14[256*13+10], codeword_reg13[256*13+10], codeword_reg12[256*13+10], codeword_reg11[256*13+10], codeword_reg10[256*13+10], codeword_reg9[256*13+10], codeword_reg8[256*13+10], codeword_reg7[256*13+10], codeword_reg6[256*13+10], codeword_reg5[256*13+10], codeword_reg4[256*13+10], codeword_reg3[256*13+10], codeword_reg2[256*13+10], codeword_reg1[256*13+10], codeword_reg16[256*12+10], codeword_reg15[256*12+10], codeword_reg14[256*12+10], codeword_reg13[256*12+10], codeword_reg12[256*12+10], codeword_reg11[256*12+10], codeword_reg10[256*12+10], codeword_reg9[256*12+10], codeword_reg8[256*12+10], codeword_reg7[256*12+10], codeword_reg6[256*12+10], codeword_reg5[256*12+10], codeword_reg4[256*12+10], codeword_reg3[256*12+10], codeword_reg2[256*12+10], codeword_reg1[256*12+10], codeword_reg16[256*11+10], codeword_reg15[256*11+10], codeword_reg14[256*11+10], codeword_reg13[256*11+10], codeword_reg12[256*11+10], codeword_reg11[256*11+10], codeword_reg10[256*11+10], codeword_reg9[256*11+10], codeword_reg8[256*11+10], codeword_reg7[256*11+10], codeword_reg6[256*11+10], codeword_reg5[256*11+10], codeword_reg4[256*11+10], codeword_reg3[256*11+10], codeword_reg2[256*11+10], codeword_reg1[256*11+10], codeword_reg16[256*10+10], codeword_reg15[256*10+10], codeword_reg14[256*10+10], codeword_reg13[256*10+10], codeword_reg12[256*10+10], codeword_reg11[256*10+10], codeword_reg10[256*10+10], codeword_reg9[256*10+10], codeword_reg8[256*10+10], codeword_reg7[256*10+10], codeword_reg6[256*10+10], codeword_reg5[256*10+10], codeword_reg4[256*10+10], codeword_reg3[256*10+10], codeword_reg2[256*10+10], codeword_reg1[256*10+10], codeword_reg16[256*9+10], codeword_reg15[256*9+10], codeword_reg14[256*9+10], codeword_reg13[256*9+10], codeword_reg12[256*9+10], codeword_reg11[256*9+10], codeword_reg10[256*9+10], codeword_reg9[256*9+10], codeword_reg8[256*9+10], codeword_reg7[256*9+10], codeword_reg6[256*9+10], codeword_reg5[256*9+10], codeword_reg4[256*9+10], codeword_reg3[256*9+10], codeword_reg2[256*9+10], codeword_reg1[256*9+10], codeword_reg16[256*8+10], codeword_reg15[256*8+10], codeword_reg14[256*8+10], codeword_reg13[256*8+10], codeword_reg12[256*8+10], codeword_reg11[256*8+10], codeword_reg10[256*8+10], codeword_reg9[256*8+10], codeword_reg8[256*8+10], codeword_reg7[256*8+10], codeword_reg6[256*8+10], codeword_reg5[256*8+10], codeword_reg4[256*8+10], codeword_reg3[256*8+10], codeword_reg2[256*8+10], codeword_reg1[256*8+10], codeword_reg16[256*7+10], codeword_reg15[256*7+10], codeword_reg14[256*7+10], codeword_reg13[256*7+10], codeword_reg12[256*7+10], codeword_reg11[256*7+10], codeword_reg10[256*7+10], codeword_reg9[256*7+10], codeword_reg8[256*7+10], codeword_reg7[256*7+10], codeword_reg6[256*7+10], codeword_reg5[256*7+10], codeword_reg4[256*7+10], codeword_reg3[256*7+10], codeword_reg2[256*7+10], codeword_reg1[256*7+10], codeword_reg16[256*6+10], codeword_reg15[256*6+10], codeword_reg14[256*6+10], codeword_reg13[256*6+10], codeword_reg12[256*6+10], codeword_reg11[256*6+10], codeword_reg10[256*6+10], codeword_reg9[256*6+10], codeword_reg8[256*6+10], codeword_reg7[256*6+10], codeword_reg6[256*6+10], codeword_reg5[256*6+10], codeword_reg4[256*6+10], codeword_reg3[256*6+10], codeword_reg2[256*6+10], codeword_reg1[256*6+10], codeword_reg16[256*5+10], codeword_reg15[256*5+10], codeword_reg14[256*5+10], codeword_reg13[256*5+10], codeword_reg12[256*5+10], codeword_reg11[256*5+10], codeword_reg10[256*5+10], codeword_reg9[256*5+10], codeword_reg8[256*5+10], codeword_reg7[256*5+10], codeword_reg6[256*5+10], codeword_reg5[256*5+10], codeword_reg4[256*5+10], codeword_reg3[256*5+10], codeword_reg2[256*5+10], codeword_reg1[256*5+10], codeword_reg16[256*4+10], codeword_reg15[256*4+10], codeword_reg14[256*4+10], codeword_reg13[256*4+10], codeword_reg12[256*4+10], codeword_reg11[256*4+10], codeword_reg10[256*4+10], codeword_reg9[256*4+10], codeword_reg8[256*4+10], codeword_reg7[256*4+10], codeword_reg6[256*4+10], codeword_reg5[256*4+10], codeword_reg4[256*4+10], codeword_reg3[256*4+10], codeword_reg2[256*4+10], codeword_reg1[256*4+10], codeword_reg16[256*3+10], codeword_reg15[256*3+10], codeword_reg14[256*3+10], codeword_reg13[256*3+10], codeword_reg12[256*3+10], codeword_reg11[256*3+10], codeword_reg10[256*3+10], codeword_reg9[256*3+10], codeword_reg8[256*3+10], codeword_reg7[256*3+10], codeword_reg6[256*3+10], codeword_reg5[256*3+10], codeword_reg4[256*3+10], codeword_reg3[256*3+10], codeword_reg2[256*3+10], codeword_reg1[256*3+10], codeword_reg16[256*2+10], codeword_reg15[256*2+10], codeword_reg14[256*2+10], codeword_reg13[256*2+10], codeword_reg12[256*2+10], codeword_reg11[256*2+10], codeword_reg10[256*2+10], codeword_reg9[256*2+10], codeword_reg8[256*2+10], codeword_reg7[256*2+10], codeword_reg6[256*2+10], codeword_reg5[256*2+10], codeword_reg4[256*2+10], codeword_reg3[256*2+10], codeword_reg2[256*2+10], codeword_reg1[256*2+10], codeword_reg16[256*1+10], codeword_reg15[256*1+10], codeword_reg14[256*1+10], codeword_reg13[256*1+10], codeword_reg12[256*1+10], codeword_reg11[256*1+10], codeword_reg10[256*1+10], codeword_reg9[256*1+10], codeword_reg8[256*1+10], codeword_reg7[256*1+10], codeword_reg6[256*1+10], codeword_reg5[256*1+10], codeword_reg4[256*1+10], codeword_reg3[256*1+10], codeword_reg2[256*1+10], codeword_reg1[256*1+10], codeword_reg16[256*0+10], codeword_reg15[256*0+10], codeword_reg14[256*0+10], codeword_reg13[256*0+10], codeword_reg12[256*0+10], codeword_reg11[256*0+10], codeword_reg10[256*0+10], codeword_reg9[256*0+10], codeword_reg8[256*0+10], codeword_reg7[256*0+10], codeword_reg6[256*0+10], codeword_reg5[256*0+10], codeword_reg4[256*0+10], codeword_reg3[256*0+10], codeword_reg2[256*0+10], codeword_reg1[256*0+10]};
                                in_bits12 <= {codeword16[11], codeword15[11], codeword14[11], codeword13[11], codeword12[11], codeword11[11], codeword10[11], codeword9[11], codeword8[11], codeword7[11], codeword6[11], codeword5[11], codeword4[11], codeword3[11], codeword2[11], codeword1[11], codeword_reg16[256*13+11], codeword_reg15[256*13+11], codeword_reg14[256*13+11], codeword_reg13[256*13+11], codeword_reg12[256*13+11], codeword_reg11[256*13+11], codeword_reg10[256*13+11], codeword_reg9[256*13+11], codeword_reg8[256*13+11], codeword_reg7[256*13+11], codeword_reg6[256*13+11], codeword_reg5[256*13+11], codeword_reg4[256*13+11], codeword_reg3[256*13+11], codeword_reg2[256*13+11], codeword_reg1[256*13+11], codeword_reg16[256*12+11], codeword_reg15[256*12+11], codeword_reg14[256*12+11], codeword_reg13[256*12+11], codeword_reg12[256*12+11], codeword_reg11[256*12+11], codeword_reg10[256*12+11], codeword_reg9[256*12+11], codeword_reg8[256*12+11], codeword_reg7[256*12+11], codeword_reg6[256*12+11], codeword_reg5[256*12+11], codeword_reg4[256*12+11], codeword_reg3[256*12+11], codeword_reg2[256*12+11], codeword_reg1[256*12+11], codeword_reg16[256*11+11], codeword_reg15[256*11+11], codeword_reg14[256*11+11], codeword_reg13[256*11+11], codeword_reg12[256*11+11], codeword_reg11[256*11+11], codeword_reg10[256*11+11], codeword_reg9[256*11+11], codeword_reg8[256*11+11], codeword_reg7[256*11+11], codeword_reg6[256*11+11], codeword_reg5[256*11+11], codeword_reg4[256*11+11], codeword_reg3[256*11+11], codeword_reg2[256*11+11], codeword_reg1[256*11+11], codeword_reg16[256*10+11], codeword_reg15[256*10+11], codeword_reg14[256*10+11], codeword_reg13[256*10+11], codeword_reg12[256*10+11], codeword_reg11[256*10+11], codeword_reg10[256*10+11], codeword_reg9[256*10+11], codeword_reg8[256*10+11], codeword_reg7[256*10+11], codeword_reg6[256*10+11], codeword_reg5[256*10+11], codeword_reg4[256*10+11], codeword_reg3[256*10+11], codeword_reg2[256*10+11], codeword_reg1[256*10+11], codeword_reg16[256*9+11], codeword_reg15[256*9+11], codeword_reg14[256*9+11], codeword_reg13[256*9+11], codeword_reg12[256*9+11], codeword_reg11[256*9+11], codeword_reg10[256*9+11], codeword_reg9[256*9+11], codeword_reg8[256*9+11], codeword_reg7[256*9+11], codeword_reg6[256*9+11], codeword_reg5[256*9+11], codeword_reg4[256*9+11], codeword_reg3[256*9+11], codeword_reg2[256*9+11], codeword_reg1[256*9+11], codeword_reg16[256*8+11], codeword_reg15[256*8+11], codeword_reg14[256*8+11], codeword_reg13[256*8+11], codeword_reg12[256*8+11], codeword_reg11[256*8+11], codeword_reg10[256*8+11], codeword_reg9[256*8+11], codeword_reg8[256*8+11], codeword_reg7[256*8+11], codeword_reg6[256*8+11], codeword_reg5[256*8+11], codeword_reg4[256*8+11], codeword_reg3[256*8+11], codeword_reg2[256*8+11], codeword_reg1[256*8+11], codeword_reg16[256*7+11], codeword_reg15[256*7+11], codeword_reg14[256*7+11], codeword_reg13[256*7+11], codeword_reg12[256*7+11], codeword_reg11[256*7+11], codeword_reg10[256*7+11], codeword_reg9[256*7+11], codeword_reg8[256*7+11], codeword_reg7[256*7+11], codeword_reg6[256*7+11], codeword_reg5[256*7+11], codeword_reg4[256*7+11], codeword_reg3[256*7+11], codeword_reg2[256*7+11], codeword_reg1[256*7+11], codeword_reg16[256*6+11], codeword_reg15[256*6+11], codeword_reg14[256*6+11], codeword_reg13[256*6+11], codeword_reg12[256*6+11], codeword_reg11[256*6+11], codeword_reg10[256*6+11], codeword_reg9[256*6+11], codeword_reg8[256*6+11], codeword_reg7[256*6+11], codeword_reg6[256*6+11], codeword_reg5[256*6+11], codeword_reg4[256*6+11], codeword_reg3[256*6+11], codeword_reg2[256*6+11], codeword_reg1[256*6+11], codeword_reg16[256*5+11], codeword_reg15[256*5+11], codeword_reg14[256*5+11], codeword_reg13[256*5+11], codeword_reg12[256*5+11], codeword_reg11[256*5+11], codeword_reg10[256*5+11], codeword_reg9[256*5+11], codeword_reg8[256*5+11], codeword_reg7[256*5+11], codeword_reg6[256*5+11], codeword_reg5[256*5+11], codeword_reg4[256*5+11], codeword_reg3[256*5+11], codeword_reg2[256*5+11], codeword_reg1[256*5+11], codeword_reg16[256*4+11], codeword_reg15[256*4+11], codeword_reg14[256*4+11], codeword_reg13[256*4+11], codeword_reg12[256*4+11], codeword_reg11[256*4+11], codeword_reg10[256*4+11], codeword_reg9[256*4+11], codeword_reg8[256*4+11], codeword_reg7[256*4+11], codeword_reg6[256*4+11], codeword_reg5[256*4+11], codeword_reg4[256*4+11], codeword_reg3[256*4+11], codeword_reg2[256*4+11], codeword_reg1[256*4+11], codeword_reg16[256*3+11], codeword_reg15[256*3+11], codeword_reg14[256*3+11], codeword_reg13[256*3+11], codeword_reg12[256*3+11], codeword_reg11[256*3+11], codeword_reg10[256*3+11], codeword_reg9[256*3+11], codeword_reg8[256*3+11], codeword_reg7[256*3+11], codeword_reg6[256*3+11], codeword_reg5[256*3+11], codeword_reg4[256*3+11], codeword_reg3[256*3+11], codeword_reg2[256*3+11], codeword_reg1[256*3+11], codeword_reg16[256*2+11], codeword_reg15[256*2+11], codeword_reg14[256*2+11], codeword_reg13[256*2+11], codeword_reg12[256*2+11], codeword_reg11[256*2+11], codeword_reg10[256*2+11], codeword_reg9[256*2+11], codeword_reg8[256*2+11], codeword_reg7[256*2+11], codeword_reg6[256*2+11], codeword_reg5[256*2+11], codeword_reg4[256*2+11], codeword_reg3[256*2+11], codeword_reg2[256*2+11], codeword_reg1[256*2+11], codeword_reg16[256*1+11], codeword_reg15[256*1+11], codeword_reg14[256*1+11], codeword_reg13[256*1+11], codeword_reg12[256*1+11], codeword_reg11[256*1+11], codeword_reg10[256*1+11], codeword_reg9[256*1+11], codeword_reg8[256*1+11], codeword_reg7[256*1+11], codeword_reg6[256*1+11], codeword_reg5[256*1+11], codeword_reg4[256*1+11], codeword_reg3[256*1+11], codeword_reg2[256*1+11], codeword_reg1[256*1+11], codeword_reg16[256*0+11], codeword_reg15[256*0+11], codeword_reg14[256*0+11], codeword_reg13[256*0+11], codeword_reg12[256*0+11], codeword_reg11[256*0+11], codeword_reg10[256*0+11], codeword_reg9[256*0+11], codeword_reg8[256*0+11], codeword_reg7[256*0+11], codeword_reg6[256*0+11], codeword_reg5[256*0+11], codeword_reg4[256*0+11], codeword_reg3[256*0+11], codeword_reg2[256*0+11], codeword_reg1[256*0+11]};
                                in_bits13 <= {codeword16[12], codeword15[12], codeword14[12], codeword13[12], codeword12[12], codeword11[12], codeword10[12], codeword9[12], codeword8[12], codeword7[12], codeword6[12], codeword5[12], codeword4[12], codeword3[12], codeword2[12], codeword1[12], codeword_reg16[256*13+12], codeword_reg15[256*13+12], codeword_reg14[256*13+12], codeword_reg13[256*13+12], codeword_reg12[256*13+12], codeword_reg11[256*13+12], codeword_reg10[256*13+12], codeword_reg9[256*13+12], codeword_reg8[256*13+12], codeword_reg7[256*13+12], codeword_reg6[256*13+12], codeword_reg5[256*13+12], codeword_reg4[256*13+12], codeword_reg3[256*13+12], codeword_reg2[256*13+12], codeword_reg1[256*13+12], codeword_reg16[256*12+12], codeword_reg15[256*12+12], codeword_reg14[256*12+12], codeword_reg13[256*12+12], codeword_reg12[256*12+12], codeword_reg11[256*12+12], codeword_reg10[256*12+12], codeword_reg9[256*12+12], codeword_reg8[256*12+12], codeword_reg7[256*12+12], codeword_reg6[256*12+12], codeword_reg5[256*12+12], codeword_reg4[256*12+12], codeword_reg3[256*12+12], codeword_reg2[256*12+12], codeword_reg1[256*12+12], codeword_reg16[256*11+12], codeword_reg15[256*11+12], codeword_reg14[256*11+12], codeword_reg13[256*11+12], codeword_reg12[256*11+12], codeword_reg11[256*11+12], codeword_reg10[256*11+12], codeword_reg9[256*11+12], codeword_reg8[256*11+12], codeword_reg7[256*11+12], codeword_reg6[256*11+12], codeword_reg5[256*11+12], codeword_reg4[256*11+12], codeword_reg3[256*11+12], codeword_reg2[256*11+12], codeword_reg1[256*11+12], codeword_reg16[256*10+12], codeword_reg15[256*10+12], codeword_reg14[256*10+12], codeword_reg13[256*10+12], codeword_reg12[256*10+12], codeword_reg11[256*10+12], codeword_reg10[256*10+12], codeword_reg9[256*10+12], codeword_reg8[256*10+12], codeword_reg7[256*10+12], codeword_reg6[256*10+12], codeword_reg5[256*10+12], codeword_reg4[256*10+12], codeword_reg3[256*10+12], codeword_reg2[256*10+12], codeword_reg1[256*10+12], codeword_reg16[256*9+12], codeword_reg15[256*9+12], codeword_reg14[256*9+12], codeword_reg13[256*9+12], codeword_reg12[256*9+12], codeword_reg11[256*9+12], codeword_reg10[256*9+12], codeword_reg9[256*9+12], codeword_reg8[256*9+12], codeword_reg7[256*9+12], codeword_reg6[256*9+12], codeword_reg5[256*9+12], codeword_reg4[256*9+12], codeword_reg3[256*9+12], codeword_reg2[256*9+12], codeword_reg1[256*9+12], codeword_reg16[256*8+12], codeword_reg15[256*8+12], codeword_reg14[256*8+12], codeword_reg13[256*8+12], codeword_reg12[256*8+12], codeword_reg11[256*8+12], codeword_reg10[256*8+12], codeword_reg9[256*8+12], codeword_reg8[256*8+12], codeword_reg7[256*8+12], codeword_reg6[256*8+12], codeword_reg5[256*8+12], codeword_reg4[256*8+12], codeword_reg3[256*8+12], codeword_reg2[256*8+12], codeword_reg1[256*8+12], codeword_reg16[256*7+12], codeword_reg15[256*7+12], codeword_reg14[256*7+12], codeword_reg13[256*7+12], codeword_reg12[256*7+12], codeword_reg11[256*7+12], codeword_reg10[256*7+12], codeword_reg9[256*7+12], codeword_reg8[256*7+12], codeword_reg7[256*7+12], codeword_reg6[256*7+12], codeword_reg5[256*7+12], codeword_reg4[256*7+12], codeword_reg3[256*7+12], codeword_reg2[256*7+12], codeword_reg1[256*7+12], codeword_reg16[256*6+12], codeword_reg15[256*6+12], codeword_reg14[256*6+12], codeword_reg13[256*6+12], codeword_reg12[256*6+12], codeword_reg11[256*6+12], codeword_reg10[256*6+12], codeword_reg9[256*6+12], codeword_reg8[256*6+12], codeword_reg7[256*6+12], codeword_reg6[256*6+12], codeword_reg5[256*6+12], codeword_reg4[256*6+12], codeword_reg3[256*6+12], codeword_reg2[256*6+12], codeword_reg1[256*6+12], codeword_reg16[256*5+12], codeword_reg15[256*5+12], codeword_reg14[256*5+12], codeword_reg13[256*5+12], codeword_reg12[256*5+12], codeword_reg11[256*5+12], codeword_reg10[256*5+12], codeword_reg9[256*5+12], codeword_reg8[256*5+12], codeword_reg7[256*5+12], codeword_reg6[256*5+12], codeword_reg5[256*5+12], codeword_reg4[256*5+12], codeword_reg3[256*5+12], codeword_reg2[256*5+12], codeword_reg1[256*5+12], codeword_reg16[256*4+12], codeword_reg15[256*4+12], codeword_reg14[256*4+12], codeword_reg13[256*4+12], codeword_reg12[256*4+12], codeword_reg11[256*4+12], codeword_reg10[256*4+12], codeword_reg9[256*4+12], codeword_reg8[256*4+12], codeword_reg7[256*4+12], codeword_reg6[256*4+12], codeword_reg5[256*4+12], codeword_reg4[256*4+12], codeword_reg3[256*4+12], codeword_reg2[256*4+12], codeword_reg1[256*4+12], codeword_reg16[256*3+12], codeword_reg15[256*3+12], codeword_reg14[256*3+12], codeword_reg13[256*3+12], codeword_reg12[256*3+12], codeword_reg11[256*3+12], codeword_reg10[256*3+12], codeword_reg9[256*3+12], codeword_reg8[256*3+12], codeword_reg7[256*3+12], codeword_reg6[256*3+12], codeword_reg5[256*3+12], codeword_reg4[256*3+12], codeword_reg3[256*3+12], codeword_reg2[256*3+12], codeword_reg1[256*3+12], codeword_reg16[256*2+12], codeword_reg15[256*2+12], codeword_reg14[256*2+12], codeword_reg13[256*2+12], codeword_reg12[256*2+12], codeword_reg11[256*2+12], codeword_reg10[256*2+12], codeword_reg9[256*2+12], codeword_reg8[256*2+12], codeword_reg7[256*2+12], codeword_reg6[256*2+12], codeword_reg5[256*2+12], codeword_reg4[256*2+12], codeword_reg3[256*2+12], codeword_reg2[256*2+12], codeword_reg1[256*2+12], codeword_reg16[256*1+12], codeword_reg15[256*1+12], codeword_reg14[256*1+12], codeword_reg13[256*1+12], codeword_reg12[256*1+12], codeword_reg11[256*1+12], codeword_reg10[256*1+12], codeword_reg9[256*1+12], codeword_reg8[256*1+12], codeword_reg7[256*1+12], codeword_reg6[256*1+12], codeword_reg5[256*1+12], codeword_reg4[256*1+12], codeword_reg3[256*1+12], codeword_reg2[256*1+12], codeword_reg1[256*1+12], codeword_reg16[256*0+12], codeword_reg15[256*0+12], codeword_reg14[256*0+12], codeword_reg13[256*0+12], codeword_reg12[256*0+12], codeword_reg11[256*0+12], codeword_reg10[256*0+12], codeword_reg9[256*0+12], codeword_reg8[256*0+12], codeword_reg7[256*0+12], codeword_reg6[256*0+12], codeword_reg5[256*0+12], codeword_reg4[256*0+12], codeword_reg3[256*0+12], codeword_reg2[256*0+12], codeword_reg1[256*0+12]};
                                in_bits14 <= {codeword16[13], codeword15[13], codeword14[13], codeword13[13], codeword12[13], codeword11[13], codeword10[13], codeword9[13], codeword8[13], codeword7[13], codeword6[13], codeword5[13], codeword4[13], codeword3[13], codeword2[13], codeword1[13], codeword_reg16[256*13+13], codeword_reg15[256*13+13], codeword_reg14[256*13+13], codeword_reg13[256*13+13], codeword_reg12[256*13+13], codeword_reg11[256*13+13], codeword_reg10[256*13+13], codeword_reg9[256*13+13], codeword_reg8[256*13+13], codeword_reg7[256*13+13], codeword_reg6[256*13+13], codeword_reg5[256*13+13], codeword_reg4[256*13+13], codeword_reg3[256*13+13], codeword_reg2[256*13+13], codeword_reg1[256*13+13], codeword_reg16[256*12+13], codeword_reg15[256*12+13], codeword_reg14[256*12+13], codeword_reg13[256*12+13], codeword_reg12[256*12+13], codeword_reg11[256*12+13], codeword_reg10[256*12+13], codeword_reg9[256*12+13], codeword_reg8[256*12+13], codeword_reg7[256*12+13], codeword_reg6[256*12+13], codeword_reg5[256*12+13], codeword_reg4[256*12+13], codeword_reg3[256*12+13], codeword_reg2[256*12+13], codeword_reg1[256*12+13], codeword_reg16[256*11+13], codeword_reg15[256*11+13], codeword_reg14[256*11+13], codeword_reg13[256*11+13], codeword_reg12[256*11+13], codeword_reg11[256*11+13], codeword_reg10[256*11+13], codeword_reg9[256*11+13], codeword_reg8[256*11+13], codeword_reg7[256*11+13], codeword_reg6[256*11+13], codeword_reg5[256*11+13], codeword_reg4[256*11+13], codeword_reg3[256*11+13], codeword_reg2[256*11+13], codeword_reg1[256*11+13], codeword_reg16[256*10+13], codeword_reg15[256*10+13], codeword_reg14[256*10+13], codeword_reg13[256*10+13], codeword_reg12[256*10+13], codeword_reg11[256*10+13], codeword_reg10[256*10+13], codeword_reg9[256*10+13], codeword_reg8[256*10+13], codeword_reg7[256*10+13], codeword_reg6[256*10+13], codeword_reg5[256*10+13], codeword_reg4[256*10+13], codeword_reg3[256*10+13], codeword_reg2[256*10+13], codeword_reg1[256*10+13], codeword_reg16[256*9+13], codeword_reg15[256*9+13], codeword_reg14[256*9+13], codeword_reg13[256*9+13], codeword_reg12[256*9+13], codeword_reg11[256*9+13], codeword_reg10[256*9+13], codeword_reg9[256*9+13], codeword_reg8[256*9+13], codeword_reg7[256*9+13], codeword_reg6[256*9+13], codeword_reg5[256*9+13], codeword_reg4[256*9+13], codeword_reg3[256*9+13], codeword_reg2[256*9+13], codeword_reg1[256*9+13], codeword_reg16[256*8+13], codeword_reg15[256*8+13], codeword_reg14[256*8+13], codeword_reg13[256*8+13], codeword_reg12[256*8+13], codeword_reg11[256*8+13], codeword_reg10[256*8+13], codeword_reg9[256*8+13], codeword_reg8[256*8+13], codeword_reg7[256*8+13], codeword_reg6[256*8+13], codeword_reg5[256*8+13], codeword_reg4[256*8+13], codeword_reg3[256*8+13], codeword_reg2[256*8+13], codeword_reg1[256*8+13], codeword_reg16[256*7+13], codeword_reg15[256*7+13], codeword_reg14[256*7+13], codeword_reg13[256*7+13], codeword_reg12[256*7+13], codeword_reg11[256*7+13], codeword_reg10[256*7+13], codeword_reg9[256*7+13], codeword_reg8[256*7+13], codeword_reg7[256*7+13], codeword_reg6[256*7+13], codeword_reg5[256*7+13], codeword_reg4[256*7+13], codeword_reg3[256*7+13], codeword_reg2[256*7+13], codeword_reg1[256*7+13], codeword_reg16[256*6+13], codeword_reg15[256*6+13], codeword_reg14[256*6+13], codeword_reg13[256*6+13], codeword_reg12[256*6+13], codeword_reg11[256*6+13], codeword_reg10[256*6+13], codeword_reg9[256*6+13], codeword_reg8[256*6+13], codeword_reg7[256*6+13], codeword_reg6[256*6+13], codeword_reg5[256*6+13], codeword_reg4[256*6+13], codeword_reg3[256*6+13], codeword_reg2[256*6+13], codeword_reg1[256*6+13], codeword_reg16[256*5+13], codeword_reg15[256*5+13], codeword_reg14[256*5+13], codeword_reg13[256*5+13], codeword_reg12[256*5+13], codeword_reg11[256*5+13], codeword_reg10[256*5+13], codeword_reg9[256*5+13], codeword_reg8[256*5+13], codeword_reg7[256*5+13], codeword_reg6[256*5+13], codeword_reg5[256*5+13], codeword_reg4[256*5+13], codeword_reg3[256*5+13], codeword_reg2[256*5+13], codeword_reg1[256*5+13], codeword_reg16[256*4+13], codeword_reg15[256*4+13], codeword_reg14[256*4+13], codeword_reg13[256*4+13], codeword_reg12[256*4+13], codeword_reg11[256*4+13], codeword_reg10[256*4+13], codeword_reg9[256*4+13], codeword_reg8[256*4+13], codeword_reg7[256*4+13], codeword_reg6[256*4+13], codeword_reg5[256*4+13], codeword_reg4[256*4+13], codeword_reg3[256*4+13], codeword_reg2[256*4+13], codeword_reg1[256*4+13], codeword_reg16[256*3+13], codeword_reg15[256*3+13], codeword_reg14[256*3+13], codeword_reg13[256*3+13], codeword_reg12[256*3+13], codeword_reg11[256*3+13], codeword_reg10[256*3+13], codeword_reg9[256*3+13], codeword_reg8[256*3+13], codeword_reg7[256*3+13], codeword_reg6[256*3+13], codeword_reg5[256*3+13], codeword_reg4[256*3+13], codeword_reg3[256*3+13], codeword_reg2[256*3+13], codeword_reg1[256*3+13], codeword_reg16[256*2+13], codeword_reg15[256*2+13], codeword_reg14[256*2+13], codeword_reg13[256*2+13], codeword_reg12[256*2+13], codeword_reg11[256*2+13], codeword_reg10[256*2+13], codeword_reg9[256*2+13], codeword_reg8[256*2+13], codeword_reg7[256*2+13], codeword_reg6[256*2+13], codeword_reg5[256*2+13], codeword_reg4[256*2+13], codeword_reg3[256*2+13], codeword_reg2[256*2+13], codeword_reg1[256*2+13], codeword_reg16[256*1+13], codeword_reg15[256*1+13], codeword_reg14[256*1+13], codeword_reg13[256*1+13], codeword_reg12[256*1+13], codeword_reg11[256*1+13], codeword_reg10[256*1+13], codeword_reg9[256*1+13], codeword_reg8[256*1+13], codeword_reg7[256*1+13], codeword_reg6[256*1+13], codeword_reg5[256*1+13], codeword_reg4[256*1+13], codeword_reg3[256*1+13], codeword_reg2[256*1+13], codeword_reg1[256*1+13], codeword_reg16[256*0+13], codeword_reg15[256*0+13], codeword_reg14[256*0+13], codeword_reg13[256*0+13], codeword_reg12[256*0+13], codeword_reg11[256*0+13], codeword_reg10[256*0+13], codeword_reg9[256*0+13], codeword_reg8[256*0+13], codeword_reg7[256*0+13], codeword_reg6[256*0+13], codeword_reg5[256*0+13], codeword_reg4[256*0+13], codeword_reg3[256*0+13], codeword_reg2[256*0+13], codeword_reg1[256*0+13]};
                                in_bits15 <= {codeword16[14], codeword15[14], codeword14[14], codeword13[14], codeword12[14], codeword11[14], codeword10[14], codeword9[14], codeword8[14], codeword7[14], codeword6[14], codeword5[14], codeword4[14], codeword3[14], codeword2[14], codeword1[14], codeword_reg16[256*13+14], codeword_reg15[256*13+14], codeword_reg14[256*13+14], codeword_reg13[256*13+14], codeword_reg12[256*13+14], codeword_reg11[256*13+14], codeword_reg10[256*13+14], codeword_reg9[256*13+14], codeword_reg8[256*13+14], codeword_reg7[256*13+14], codeword_reg6[256*13+14], codeword_reg5[256*13+14], codeword_reg4[256*13+14], codeword_reg3[256*13+14], codeword_reg2[256*13+14], codeword_reg1[256*13+14], codeword_reg16[256*12+14], codeword_reg15[256*12+14], codeword_reg14[256*12+14], codeword_reg13[256*12+14], codeword_reg12[256*12+14], codeword_reg11[256*12+14], codeword_reg10[256*12+14], codeword_reg9[256*12+14], codeword_reg8[256*12+14], codeword_reg7[256*12+14], codeword_reg6[256*12+14], codeword_reg5[256*12+14], codeword_reg4[256*12+14], codeword_reg3[256*12+14], codeword_reg2[256*12+14], codeword_reg1[256*12+14], codeword_reg16[256*11+14], codeword_reg15[256*11+14], codeword_reg14[256*11+14], codeword_reg13[256*11+14], codeword_reg12[256*11+14], codeword_reg11[256*11+14], codeword_reg10[256*11+14], codeword_reg9[256*11+14], codeword_reg8[256*11+14], codeword_reg7[256*11+14], codeword_reg6[256*11+14], codeword_reg5[256*11+14], codeword_reg4[256*11+14], codeword_reg3[256*11+14], codeword_reg2[256*11+14], codeword_reg1[256*11+14], codeword_reg16[256*10+14], codeword_reg15[256*10+14], codeword_reg14[256*10+14], codeword_reg13[256*10+14], codeword_reg12[256*10+14], codeword_reg11[256*10+14], codeword_reg10[256*10+14], codeword_reg9[256*10+14], codeword_reg8[256*10+14], codeword_reg7[256*10+14], codeword_reg6[256*10+14], codeword_reg5[256*10+14], codeword_reg4[256*10+14], codeword_reg3[256*10+14], codeword_reg2[256*10+14], codeword_reg1[256*10+14], codeword_reg16[256*9+14], codeword_reg15[256*9+14], codeword_reg14[256*9+14], codeword_reg13[256*9+14], codeword_reg12[256*9+14], codeword_reg11[256*9+14], codeword_reg10[256*9+14], codeword_reg9[256*9+14], codeword_reg8[256*9+14], codeword_reg7[256*9+14], codeword_reg6[256*9+14], codeword_reg5[256*9+14], codeword_reg4[256*9+14], codeword_reg3[256*9+14], codeword_reg2[256*9+14], codeword_reg1[256*9+14], codeword_reg16[256*8+14], codeword_reg15[256*8+14], codeword_reg14[256*8+14], codeword_reg13[256*8+14], codeword_reg12[256*8+14], codeword_reg11[256*8+14], codeword_reg10[256*8+14], codeword_reg9[256*8+14], codeword_reg8[256*8+14], codeword_reg7[256*8+14], codeword_reg6[256*8+14], codeword_reg5[256*8+14], codeword_reg4[256*8+14], codeword_reg3[256*8+14], codeword_reg2[256*8+14], codeword_reg1[256*8+14], codeword_reg16[256*7+14], codeword_reg15[256*7+14], codeword_reg14[256*7+14], codeword_reg13[256*7+14], codeword_reg12[256*7+14], codeword_reg11[256*7+14], codeword_reg10[256*7+14], codeword_reg9[256*7+14], codeword_reg8[256*7+14], codeword_reg7[256*7+14], codeword_reg6[256*7+14], codeword_reg5[256*7+14], codeword_reg4[256*7+14], codeword_reg3[256*7+14], codeword_reg2[256*7+14], codeword_reg1[256*7+14], codeword_reg16[256*6+14], codeword_reg15[256*6+14], codeword_reg14[256*6+14], codeword_reg13[256*6+14], codeword_reg12[256*6+14], codeword_reg11[256*6+14], codeword_reg10[256*6+14], codeword_reg9[256*6+14], codeword_reg8[256*6+14], codeword_reg7[256*6+14], codeword_reg6[256*6+14], codeword_reg5[256*6+14], codeword_reg4[256*6+14], codeword_reg3[256*6+14], codeword_reg2[256*6+14], codeword_reg1[256*6+14], codeword_reg16[256*5+14], codeword_reg15[256*5+14], codeword_reg14[256*5+14], codeword_reg13[256*5+14], codeword_reg12[256*5+14], codeword_reg11[256*5+14], codeword_reg10[256*5+14], codeword_reg9[256*5+14], codeword_reg8[256*5+14], codeword_reg7[256*5+14], codeword_reg6[256*5+14], codeword_reg5[256*5+14], codeword_reg4[256*5+14], codeword_reg3[256*5+14], codeword_reg2[256*5+14], codeword_reg1[256*5+14], codeword_reg16[256*4+14], codeword_reg15[256*4+14], codeword_reg14[256*4+14], codeword_reg13[256*4+14], codeword_reg12[256*4+14], codeword_reg11[256*4+14], codeword_reg10[256*4+14], codeword_reg9[256*4+14], codeword_reg8[256*4+14], codeword_reg7[256*4+14], codeword_reg6[256*4+14], codeword_reg5[256*4+14], codeword_reg4[256*4+14], codeword_reg3[256*4+14], codeword_reg2[256*4+14], codeword_reg1[256*4+14], codeword_reg16[256*3+14], codeword_reg15[256*3+14], codeword_reg14[256*3+14], codeword_reg13[256*3+14], codeword_reg12[256*3+14], codeword_reg11[256*3+14], codeword_reg10[256*3+14], codeword_reg9[256*3+14], codeword_reg8[256*3+14], codeword_reg7[256*3+14], codeword_reg6[256*3+14], codeword_reg5[256*3+14], codeword_reg4[256*3+14], codeword_reg3[256*3+14], codeword_reg2[256*3+14], codeword_reg1[256*3+14], codeword_reg16[256*2+14], codeword_reg15[256*2+14], codeword_reg14[256*2+14], codeword_reg13[256*2+14], codeword_reg12[256*2+14], codeword_reg11[256*2+14], codeword_reg10[256*2+14], codeword_reg9[256*2+14], codeword_reg8[256*2+14], codeword_reg7[256*2+14], codeword_reg6[256*2+14], codeword_reg5[256*2+14], codeword_reg4[256*2+14], codeword_reg3[256*2+14], codeword_reg2[256*2+14], codeword_reg1[256*2+14], codeword_reg16[256*1+14], codeword_reg15[256*1+14], codeword_reg14[256*1+14], codeword_reg13[256*1+14], codeword_reg12[256*1+14], codeword_reg11[256*1+14], codeword_reg10[256*1+14], codeword_reg9[256*1+14], codeword_reg8[256*1+14], codeword_reg7[256*1+14], codeword_reg6[256*1+14], codeword_reg5[256*1+14], codeword_reg4[256*1+14], codeword_reg3[256*1+14], codeword_reg2[256*1+14], codeword_reg1[256*1+14], codeword_reg16[256*0+14], codeword_reg15[256*0+14], codeword_reg14[256*0+14], codeword_reg13[256*0+14], codeword_reg12[256*0+14], codeword_reg11[256*0+14], codeword_reg10[256*0+14], codeword_reg9[256*0+14], codeword_reg8[256*0+14], codeword_reg7[256*0+14], codeword_reg6[256*0+14], codeword_reg5[256*0+14], codeword_reg4[256*0+14], codeword_reg3[256*0+14], codeword_reg2[256*0+14], codeword_reg1[256*0+14]};
                                in_bits16 <= {codeword16[15], codeword15[15], codeword14[15], codeword13[15], codeword12[15], codeword11[15], codeword10[15], codeword9[15], codeword8[15], codeword7[15], codeword6[15], codeword5[15], codeword4[15], codeword3[15], codeword2[15], codeword1[15], codeword_reg16[256*13+15], codeword_reg15[256*13+15], codeword_reg14[256*13+15], codeword_reg13[256*13+15], codeword_reg12[256*13+15], codeword_reg11[256*13+15], codeword_reg10[256*13+15], codeword_reg9[256*13+15], codeword_reg8[256*13+15], codeword_reg7[256*13+15], codeword_reg6[256*13+15], codeword_reg5[256*13+15], codeword_reg4[256*13+15], codeword_reg3[256*13+15], codeword_reg2[256*13+15], codeword_reg1[256*13+15], codeword_reg16[256*12+15], codeword_reg15[256*12+15], codeword_reg14[256*12+15], codeword_reg13[256*12+15], codeword_reg12[256*12+15], codeword_reg11[256*12+15], codeword_reg10[256*12+15], codeword_reg9[256*12+15], codeword_reg8[256*12+15], codeword_reg7[256*12+15], codeword_reg6[256*12+15], codeword_reg5[256*12+15], codeword_reg4[256*12+15], codeword_reg3[256*12+15], codeword_reg2[256*12+15], codeword_reg1[256*12+15], codeword_reg16[256*11+15], codeword_reg15[256*11+15], codeword_reg14[256*11+15], codeword_reg13[256*11+15], codeword_reg12[256*11+15], codeword_reg11[256*11+15], codeword_reg10[256*11+15], codeword_reg9[256*11+15], codeword_reg8[256*11+15], codeword_reg7[256*11+15], codeword_reg6[256*11+15], codeword_reg5[256*11+15], codeword_reg4[256*11+15], codeword_reg3[256*11+15], codeword_reg2[256*11+15], codeword_reg1[256*11+15], codeword_reg16[256*10+15], codeword_reg15[256*10+15], codeword_reg14[256*10+15], codeword_reg13[256*10+15], codeword_reg12[256*10+15], codeword_reg11[256*10+15], codeword_reg10[256*10+15], codeword_reg9[256*10+15], codeword_reg8[256*10+15], codeword_reg7[256*10+15], codeword_reg6[256*10+15], codeword_reg5[256*10+15], codeword_reg4[256*10+15], codeword_reg3[256*10+15], codeword_reg2[256*10+15], codeword_reg1[256*10+15], codeword_reg16[256*9+15], codeword_reg15[256*9+15], codeword_reg14[256*9+15], codeword_reg13[256*9+15], codeword_reg12[256*9+15], codeword_reg11[256*9+15], codeword_reg10[256*9+15], codeword_reg9[256*9+15], codeword_reg8[256*9+15], codeword_reg7[256*9+15], codeword_reg6[256*9+15], codeword_reg5[256*9+15], codeword_reg4[256*9+15], codeword_reg3[256*9+15], codeword_reg2[256*9+15], codeword_reg1[256*9+15], codeword_reg16[256*8+15], codeword_reg15[256*8+15], codeword_reg14[256*8+15], codeword_reg13[256*8+15], codeword_reg12[256*8+15], codeword_reg11[256*8+15], codeword_reg10[256*8+15], codeword_reg9[256*8+15], codeword_reg8[256*8+15], codeword_reg7[256*8+15], codeword_reg6[256*8+15], codeword_reg5[256*8+15], codeword_reg4[256*8+15], codeword_reg3[256*8+15], codeword_reg2[256*8+15], codeword_reg1[256*8+15], codeword_reg16[256*7+15], codeword_reg15[256*7+15], codeword_reg14[256*7+15], codeword_reg13[256*7+15], codeword_reg12[256*7+15], codeword_reg11[256*7+15], codeword_reg10[256*7+15], codeword_reg9[256*7+15], codeword_reg8[256*7+15], codeword_reg7[256*7+15], codeword_reg6[256*7+15], codeword_reg5[256*7+15], codeword_reg4[256*7+15], codeword_reg3[256*7+15], codeword_reg2[256*7+15], codeword_reg1[256*7+15], codeword_reg16[256*6+15], codeword_reg15[256*6+15], codeword_reg14[256*6+15], codeword_reg13[256*6+15], codeword_reg12[256*6+15], codeword_reg11[256*6+15], codeword_reg10[256*6+15], codeword_reg9[256*6+15], codeword_reg8[256*6+15], codeword_reg7[256*6+15], codeword_reg6[256*6+15], codeword_reg5[256*6+15], codeword_reg4[256*6+15], codeword_reg3[256*6+15], codeword_reg2[256*6+15], codeword_reg1[256*6+15], codeword_reg16[256*5+15], codeword_reg15[256*5+15], codeword_reg14[256*5+15], codeword_reg13[256*5+15], codeword_reg12[256*5+15], codeword_reg11[256*5+15], codeword_reg10[256*5+15], codeword_reg9[256*5+15], codeword_reg8[256*5+15], codeword_reg7[256*5+15], codeword_reg6[256*5+15], codeword_reg5[256*5+15], codeword_reg4[256*5+15], codeword_reg3[256*5+15], codeword_reg2[256*5+15], codeword_reg1[256*5+15], codeword_reg16[256*4+15], codeword_reg15[256*4+15], codeword_reg14[256*4+15], codeword_reg13[256*4+15], codeword_reg12[256*4+15], codeword_reg11[256*4+15], codeword_reg10[256*4+15], codeword_reg9[256*4+15], codeword_reg8[256*4+15], codeword_reg7[256*4+15], codeword_reg6[256*4+15], codeword_reg5[256*4+15], codeword_reg4[256*4+15], codeword_reg3[256*4+15], codeword_reg2[256*4+15], codeword_reg1[256*4+15], codeword_reg16[256*3+15], codeword_reg15[256*3+15], codeword_reg14[256*3+15], codeword_reg13[256*3+15], codeword_reg12[256*3+15], codeword_reg11[256*3+15], codeword_reg10[256*3+15], codeword_reg9[256*3+15], codeword_reg8[256*3+15], codeword_reg7[256*3+15], codeword_reg6[256*3+15], codeword_reg5[256*3+15], codeword_reg4[256*3+15], codeword_reg3[256*3+15], codeword_reg2[256*3+15], codeword_reg1[256*3+15], codeword_reg16[256*2+15], codeword_reg15[256*2+15], codeword_reg14[256*2+15], codeword_reg13[256*2+15], codeword_reg12[256*2+15], codeword_reg11[256*2+15], codeword_reg10[256*2+15], codeword_reg9[256*2+15], codeword_reg8[256*2+15], codeword_reg7[256*2+15], codeword_reg6[256*2+15], codeword_reg5[256*2+15], codeword_reg4[256*2+15], codeword_reg3[256*2+15], codeword_reg2[256*2+15], codeword_reg1[256*2+15], codeword_reg16[256*1+15], codeword_reg15[256*1+15], codeword_reg14[256*1+15], codeword_reg13[256*1+15], codeword_reg12[256*1+15], codeword_reg11[256*1+15], codeword_reg10[256*1+15], codeword_reg9[256*1+15], codeword_reg8[256*1+15], codeword_reg7[256*1+15], codeword_reg6[256*1+15], codeword_reg5[256*1+15], codeword_reg4[256*1+15], codeword_reg3[256*1+15], codeword_reg2[256*1+15], codeword_reg1[256*1+15], codeword_reg16[256*0+15], codeword_reg15[256*0+15], codeword_reg14[256*0+15], codeword_reg13[256*0+15], codeword_reg12[256*0+15], codeword_reg11[256*0+15], codeword_reg10[256*0+15], codeword_reg9[256*0+15], codeword_reg8[256*0+15], codeword_reg7[256*0+15], codeword_reg6[256*0+15], codeword_reg5[256*0+15], codeword_reg4[256*0+15], codeword_reg3[256*0+15], codeword_reg2[256*0+15], codeword_reg1[256*0+15]};
                            
                            codeword_reg1[(set_id)*n  +: n] <= codeword1;
                            codeword_reg2[(set_id)*n  +: n] <= codeword2;
                            codeword_reg3[(set_id)*n  +: n] <= codeword3;
                            codeword_reg4[(set_id)*n  +: n] <= codeword4;
                            codeword_reg5[(set_id)*n  +: n] <= codeword5;
                            codeword_reg6[(set_id)*n  +: n] <= codeword6;
                            codeword_reg7[(set_id)*n  +: n] <= codeword7;
                            codeword_reg8[(set_id)*n  +: n] <= codeword8;
                            codeword_reg9[(set_id)*n  +: n] <= codeword9;
                            codeword_reg10[(set_id)*n +: n] <= codeword10;
                            codeword_reg11[(set_id)*n +: n] <= codeword11;
                            codeword_reg12[(set_id)*n +: n] <= codeword12;
                            codeword_reg13[(set_id)*n +: n] <= codeword13;
                            codeword_reg14[(set_id)*n +: n] <= codeword14;
                            codeword_reg15[(set_id)*n +: n] <= codeword15;
                            codeword_reg16[(set_id)*n +: n] <= codeword16;
                            
                            out_codeword1  <= 'bx;
                            out_codeword2  <= 'bx;
                            out_codeword3  <= 'bx;
                            out_codeword4  <= 'bx;
                            out_codeword5  <= 'bx;
                            out_codeword6  <= 'bx;
                            out_codeword7  <= 'bx;
                            out_codeword8  <= 'bx;
                            out_codeword9  <= 'bx;
                            out_codeword10 <= 'bx;
                            out_codeword11 <= 'bx;
                            out_codeword12 <= 'bx;
                            out_codeword13 <= 'bx;
                            out_codeword14 <= 'bx;
                            out_codeword15 <= 'bx;
                            out_codeword16 <= 'bx;
                            
                            // Update the control variables
                            set_id <= 4'b1;
                            row <= 1'b0;
                            row_counter <= 4'd0;
                            new1 <= 1'b0;
                            store <= 1'b0;
                        end
                    //// End of the row encoding ////  
                        
                        
                    //// Start of the col encoding ////
                    end else begin
                    
                        // For this range of the counter, the input is taken from the buffer
                        if (col_counter < 5'd16) begin
                            
                            // Give input from the row encoded codewords using the buffer
                            in_bits1  <= {codeword_reg16[256*14+set_id*16+0], codeword_reg15[256*14+set_id*16+0], codeword_reg14[256*14+set_id*16+0], codeword_reg13[256*14+set_id*16+0], codeword_reg12[256*14+set_id*16+0], codeword_reg11[256*14+set_id*16+0], codeword_reg10[256*14+set_id*16+0], codeword_reg9[256*14+set_id*16+0], codeword_reg8[256*14+set_id*16+0], codeword_reg7[256*14+set_id*16+0], codeword_reg6[256*14+set_id*16+0], codeword_reg5[256*14+set_id*16+0], codeword_reg4[256*14+set_id*16+0], codeword_reg3[256*14+set_id*16+0], codeword_reg2[256*14+set_id*16+0], codeword_reg1[256*14+set_id*16+0], codeword_reg16[256*13+set_id*16+0], codeword_reg15[256*13+set_id*16+0], codeword_reg14[256*13+set_id*16+0], codeword_reg13[256*13+set_id*16+0], codeword_reg12[256*13+set_id*16+0], codeword_reg11[256*13+set_id*16+0], codeword_reg10[256*13+set_id*16+0], codeword_reg9[256*13+set_id*16+0], codeword_reg8[256*13+set_id*16+0], codeword_reg7[256*13+set_id*16+0], codeword_reg6[256*13+set_id*16+0], codeword_reg5[256*13+set_id*16+0], codeword_reg4[256*13+set_id*16+0], codeword_reg3[256*13+set_id*16+0], codeword_reg2[256*13+set_id*16+0], codeword_reg1[256*13+set_id*16+0], codeword_reg16[256*12+set_id*16+0], codeword_reg15[256*12+set_id*16+0], codeword_reg14[256*12+set_id*16+0], codeword_reg13[256*12+set_id*16+0], codeword_reg12[256*12+set_id*16+0], codeword_reg11[256*12+set_id*16+0], codeword_reg10[256*12+set_id*16+0], codeword_reg9[256*12+set_id*16+0], codeword_reg8[256*12+set_id*16+0], codeword_reg7[256*12+set_id*16+0], codeword_reg6[256*12+set_id*16+0], codeword_reg5[256*12+set_id*16+0], codeword_reg4[256*12+set_id*16+0], codeword_reg3[256*12+set_id*16+0], codeword_reg2[256*12+set_id*16+0], codeword_reg1[256*12+set_id*16+0], codeword_reg16[256*11+set_id*16+0], codeword_reg15[256*11+set_id*16+0], codeword_reg14[256*11+set_id*16+0], codeword_reg13[256*11+set_id*16+0], codeword_reg12[256*11+set_id*16+0], codeword_reg11[256*11+set_id*16+0], codeword_reg10[256*11+set_id*16+0], codeword_reg9[256*11+set_id*16+0], codeword_reg8[256*11+set_id*16+0], codeword_reg7[256*11+set_id*16+0], codeword_reg6[256*11+set_id*16+0], codeword_reg5[256*11+set_id*16+0], codeword_reg4[256*11+set_id*16+0], codeword_reg3[256*11+set_id*16+0], codeword_reg2[256*11+set_id*16+0], codeword_reg1[256*11+set_id*16+0], codeword_reg16[256*10+set_id*16+0], codeword_reg15[256*10+set_id*16+0], codeword_reg14[256*10+set_id*16+0], codeword_reg13[256*10+set_id*16+0], codeword_reg12[256*10+set_id*16+0], codeword_reg11[256*10+set_id*16+0], codeword_reg10[256*10+set_id*16+0], codeword_reg9[256*10+set_id*16+0], codeword_reg8[256*10+set_id*16+0], codeword_reg7[256*10+set_id*16+0], codeword_reg6[256*10+set_id*16+0], codeword_reg5[256*10+set_id*16+0], codeword_reg4[256*10+set_id*16+0], codeword_reg3[256*10+set_id*16+0], codeword_reg2[256*10+set_id*16+0], codeword_reg1[256*10+set_id*16+0], codeword_reg16[256*9+set_id*16+0], codeword_reg15[256*9+set_id*16+0], codeword_reg14[256*9+set_id*16+0], codeword_reg13[256*9+set_id*16+0], codeword_reg12[256*9+set_id*16+0], codeword_reg11[256*9+set_id*16+0], codeword_reg10[256*9+set_id*16+0], codeword_reg9[256*9+set_id*16+0], codeword_reg8[256*9+set_id*16+0], codeword_reg7[256*9+set_id*16+0], codeword_reg6[256*9+set_id*16+0], codeword_reg5[256*9+set_id*16+0], codeword_reg4[256*9+set_id*16+0], codeword_reg3[256*9+set_id*16+0], codeword_reg2[256*9+set_id*16+0], codeword_reg1[256*9+set_id*16+0], codeword_reg16[256*8+set_id*16+0], codeword_reg15[256*8+set_id*16+0], codeword_reg14[256*8+set_id*16+0], codeword_reg13[256*8+set_id*16+0], codeword_reg12[256*8+set_id*16+0], codeword_reg11[256*8+set_id*16+0], codeword_reg10[256*8+set_id*16+0], codeword_reg9[256*8+set_id*16+0], codeword_reg8[256*8+set_id*16+0], codeword_reg7[256*8+set_id*16+0], codeword_reg6[256*8+set_id*16+0], codeword_reg5[256*8+set_id*16+0], codeword_reg4[256*8+set_id*16+0], codeword_reg3[256*8+set_id*16+0], codeword_reg2[256*8+set_id*16+0], codeword_reg1[256*8+set_id*16+0], codeword_reg16[256*7+set_id*16+0], codeword_reg15[256*7+set_id*16+0], codeword_reg14[256*7+set_id*16+0], codeword_reg13[256*7+set_id*16+0], codeword_reg12[256*7+set_id*16+0], codeword_reg11[256*7+set_id*16+0], codeword_reg10[256*7+set_id*16+0], codeword_reg9[256*7+set_id*16+0], codeword_reg8[256*7+set_id*16+0], codeword_reg7[256*7+set_id*16+0], codeword_reg6[256*7+set_id*16+0], codeword_reg5[256*7+set_id*16+0], codeword_reg4[256*7+set_id*16+0], codeword_reg3[256*7+set_id*16+0], codeword_reg2[256*7+set_id*16+0], codeword_reg1[256*7+set_id*16+0], codeword_reg16[256*6+set_id*16+0], codeword_reg15[256*6+set_id*16+0], codeword_reg14[256*6+set_id*16+0], codeword_reg13[256*6+set_id*16+0], codeword_reg12[256*6+set_id*16+0], codeword_reg11[256*6+set_id*16+0], codeword_reg10[256*6+set_id*16+0], codeword_reg9[256*6+set_id*16+0], codeword_reg8[256*6+set_id*16+0], codeword_reg7[256*6+set_id*16+0], codeword_reg6[256*6+set_id*16+0], codeword_reg5[256*6+set_id*16+0], codeword_reg4[256*6+set_id*16+0], codeword_reg3[256*6+set_id*16+0], codeword_reg2[256*6+set_id*16+0], codeword_reg1[256*6+set_id*16+0], codeword_reg16[256*5+set_id*16+0], codeword_reg15[256*5+set_id*16+0], codeword_reg14[256*5+set_id*16+0], codeword_reg13[256*5+set_id*16+0], codeword_reg12[256*5+set_id*16+0], codeword_reg11[256*5+set_id*16+0], codeword_reg10[256*5+set_id*16+0], codeword_reg9[256*5+set_id*16+0], codeword_reg8[256*5+set_id*16+0], codeword_reg7[256*5+set_id*16+0], codeword_reg6[256*5+set_id*16+0], codeword_reg5[256*5+set_id*16+0], codeword_reg4[256*5+set_id*16+0], codeword_reg3[256*5+set_id*16+0], codeword_reg2[256*5+set_id*16+0], codeword_reg1[256*5+set_id*16+0], codeword_reg16[256*4+set_id*16+0], codeword_reg15[256*4+set_id*16+0], codeword_reg14[256*4+set_id*16+0], codeword_reg13[256*4+set_id*16+0], codeword_reg12[256*4+set_id*16+0], codeword_reg11[256*4+set_id*16+0], codeword_reg10[256*4+set_id*16+0], codeword_reg9[256*4+set_id*16+0], codeword_reg8[256*4+set_id*16+0], codeword_reg7[256*4+set_id*16+0], codeword_reg6[256*4+set_id*16+0], codeword_reg5[256*4+set_id*16+0], codeword_reg4[256*4+set_id*16+0], codeword_reg3[256*4+set_id*16+0], codeword_reg2[256*4+set_id*16+0], codeword_reg1[256*4+set_id*16+0], codeword_reg16[256*3+set_id*16+0], codeword_reg15[256*3+set_id*16+0], codeword_reg14[256*3+set_id*16+0], codeword_reg13[256*3+set_id*16+0], codeword_reg12[256*3+set_id*16+0], codeword_reg11[256*3+set_id*16+0], codeword_reg10[256*3+set_id*16+0], codeword_reg9[256*3+set_id*16+0], codeword_reg8[256*3+set_id*16+0], codeword_reg7[256*3+set_id*16+0], codeword_reg6[256*3+set_id*16+0], codeword_reg5[256*3+set_id*16+0], codeword_reg4[256*3+set_id*16+0], codeword_reg3[256*3+set_id*16+0], codeword_reg2[256*3+set_id*16+0], codeword_reg1[256*3+set_id*16+0], codeword_reg16[256*2+set_id*16+0], codeword_reg15[256*2+set_id*16+0], codeword_reg14[256*2+set_id*16+0], codeword_reg13[256*2+set_id*16+0], codeword_reg12[256*2+set_id*16+0], codeword_reg11[256*2+set_id*16+0], codeword_reg10[256*2+set_id*16+0], codeword_reg9[256*2+set_id*16+0], codeword_reg8[256*2+set_id*16+0], codeword_reg7[256*2+set_id*16+0], codeword_reg6[256*2+set_id*16+0], codeword_reg5[256*2+set_id*16+0], codeword_reg4[256*2+set_id*16+0], codeword_reg3[256*2+set_id*16+0], codeword_reg2[256*2+set_id*16+0], codeword_reg1[256*2+set_id*16+0], codeword_reg16[256*1+set_id*16+0], codeword_reg15[256*1+set_id*16+0], codeword_reg14[256*1+set_id*16+0], codeword_reg13[256*1+set_id*16+0], codeword_reg12[256*1+set_id*16+0], codeword_reg11[256*1+set_id*16+0], codeword_reg10[256*1+set_id*16+0], codeword_reg9[256*1+set_id*16+0], codeword_reg8[256*1+set_id*16+0], codeword_reg7[256*1+set_id*16+0], codeword_reg6[256*1+set_id*16+0], codeword_reg5[256*1+set_id*16+0], codeword_reg4[256*1+set_id*16+0], codeword_reg3[256*1+set_id*16+0], codeword_reg2[256*1+set_id*16+0], codeword_reg1[256*1+set_id*16+0], codeword_reg16[256*0+set_id*16+0], codeword_reg15[256*0+set_id*16+0], codeword_reg14[256*0+set_id*16+0], codeword_reg13[256*0+set_id*16+0], codeword_reg12[256*0+set_id*16+0], codeword_reg11[256*0+set_id*16+0], codeword_reg10[256*0+set_id*16+0], codeword_reg9[256*0+set_id*16+0], codeword_reg8[256*0+set_id*16+0], codeword_reg7[256*0+set_id*16+0], codeword_reg6[256*0+set_id*16+0], codeword_reg5[256*0+set_id*16+0], codeword_reg4[256*0+set_id*16+0], codeword_reg3[256*0+set_id*16+0], codeword_reg2[256*0+set_id*16+0], codeword_reg1[256*0+set_id*16+0]};
                            in_bits2  <= {codeword_reg16[256*14+set_id*16+1], codeword_reg15[256*14+set_id*16+1], codeword_reg14[256*14+set_id*16+1], codeword_reg13[256*14+set_id*16+1], codeword_reg12[256*14+set_id*16+1], codeword_reg11[256*14+set_id*16+1], codeword_reg10[256*14+set_id*16+1], codeword_reg9[256*14+set_id*16+1], codeword_reg8[256*14+set_id*16+1], codeword_reg7[256*14+set_id*16+1], codeword_reg6[256*14+set_id*16+1], codeword_reg5[256*14+set_id*16+1], codeword_reg4[256*14+set_id*16+1], codeword_reg3[256*14+set_id*16+1], codeword_reg2[256*14+set_id*16+1], codeword_reg1[256*14+set_id*16+1], codeword_reg16[256*13+set_id*16+1], codeword_reg15[256*13+set_id*16+1], codeword_reg14[256*13+set_id*16+1], codeword_reg13[256*13+set_id*16+1], codeword_reg12[256*13+set_id*16+1], codeword_reg11[256*13+set_id*16+1], codeword_reg10[256*13+set_id*16+1], codeword_reg9[256*13+set_id*16+1], codeword_reg8[256*13+set_id*16+1], codeword_reg7[256*13+set_id*16+1], codeword_reg6[256*13+set_id*16+1], codeword_reg5[256*13+set_id*16+1], codeword_reg4[256*13+set_id*16+1], codeword_reg3[256*13+set_id*16+1], codeword_reg2[256*13+set_id*16+1], codeword_reg1[256*13+set_id*16+1], codeword_reg16[256*12+set_id*16+1], codeword_reg15[256*12+set_id*16+1], codeword_reg14[256*12+set_id*16+1], codeword_reg13[256*12+set_id*16+1], codeword_reg12[256*12+set_id*16+1], codeword_reg11[256*12+set_id*16+1], codeword_reg10[256*12+set_id*16+1], codeword_reg9[256*12+set_id*16+1], codeword_reg8[256*12+set_id*16+1], codeword_reg7[256*12+set_id*16+1], codeword_reg6[256*12+set_id*16+1], codeword_reg5[256*12+set_id*16+1], codeword_reg4[256*12+set_id*16+1], codeword_reg3[256*12+set_id*16+1], codeword_reg2[256*12+set_id*16+1], codeword_reg1[256*12+set_id*16+1], codeword_reg16[256*11+set_id*16+1], codeword_reg15[256*11+set_id*16+1], codeword_reg14[256*11+set_id*16+1], codeword_reg13[256*11+set_id*16+1], codeword_reg12[256*11+set_id*16+1], codeword_reg11[256*11+set_id*16+1], codeword_reg10[256*11+set_id*16+1], codeword_reg9[256*11+set_id*16+1], codeword_reg8[256*11+set_id*16+1], codeword_reg7[256*11+set_id*16+1], codeword_reg6[256*11+set_id*16+1], codeword_reg5[256*11+set_id*16+1], codeword_reg4[256*11+set_id*16+1], codeword_reg3[256*11+set_id*16+1], codeword_reg2[256*11+set_id*16+1], codeword_reg1[256*11+set_id*16+1], codeword_reg16[256*10+set_id*16+1], codeword_reg15[256*10+set_id*16+1], codeword_reg14[256*10+set_id*16+1], codeword_reg13[256*10+set_id*16+1], codeword_reg12[256*10+set_id*16+1], codeword_reg11[256*10+set_id*16+1], codeword_reg10[256*10+set_id*16+1], codeword_reg9[256*10+set_id*16+1], codeword_reg8[256*10+set_id*16+1], codeword_reg7[256*10+set_id*16+1], codeword_reg6[256*10+set_id*16+1], codeword_reg5[256*10+set_id*16+1], codeword_reg4[256*10+set_id*16+1], codeword_reg3[256*10+set_id*16+1], codeword_reg2[256*10+set_id*16+1], codeword_reg1[256*10+set_id*16+1], codeword_reg16[256*9+set_id*16+1], codeword_reg15[256*9+set_id*16+1], codeword_reg14[256*9+set_id*16+1], codeword_reg13[256*9+set_id*16+1], codeword_reg12[256*9+set_id*16+1], codeword_reg11[256*9+set_id*16+1], codeword_reg10[256*9+set_id*16+1], codeword_reg9[256*9+set_id*16+1], codeword_reg8[256*9+set_id*16+1], codeword_reg7[256*9+set_id*16+1], codeword_reg6[256*9+set_id*16+1], codeword_reg5[256*9+set_id*16+1], codeword_reg4[256*9+set_id*16+1], codeword_reg3[256*9+set_id*16+1], codeword_reg2[256*9+set_id*16+1], codeword_reg1[256*9+set_id*16+1], codeword_reg16[256*8+set_id*16+1], codeword_reg15[256*8+set_id*16+1], codeword_reg14[256*8+set_id*16+1], codeword_reg13[256*8+set_id*16+1], codeword_reg12[256*8+set_id*16+1], codeword_reg11[256*8+set_id*16+1], codeword_reg10[256*8+set_id*16+1], codeword_reg9[256*8+set_id*16+1], codeword_reg8[256*8+set_id*16+1], codeword_reg7[256*8+set_id*16+1], codeword_reg6[256*8+set_id*16+1], codeword_reg5[256*8+set_id*16+1], codeword_reg4[256*8+set_id*16+1], codeword_reg3[256*8+set_id*16+1], codeword_reg2[256*8+set_id*16+1], codeword_reg1[256*8+set_id*16+1], codeword_reg16[256*7+set_id*16+1], codeword_reg15[256*7+set_id*16+1], codeword_reg14[256*7+set_id*16+1], codeword_reg13[256*7+set_id*16+1], codeword_reg12[256*7+set_id*16+1], codeword_reg11[256*7+set_id*16+1], codeword_reg10[256*7+set_id*16+1], codeword_reg9[256*7+set_id*16+1], codeword_reg8[256*7+set_id*16+1], codeword_reg7[256*7+set_id*16+1], codeword_reg6[256*7+set_id*16+1], codeword_reg5[256*7+set_id*16+1], codeword_reg4[256*7+set_id*16+1], codeword_reg3[256*7+set_id*16+1], codeword_reg2[256*7+set_id*16+1], codeword_reg1[256*7+set_id*16+1], codeword_reg16[256*6+set_id*16+1], codeword_reg15[256*6+set_id*16+1], codeword_reg14[256*6+set_id*16+1], codeword_reg13[256*6+set_id*16+1], codeword_reg12[256*6+set_id*16+1], codeword_reg11[256*6+set_id*16+1], codeword_reg10[256*6+set_id*16+1], codeword_reg9[256*6+set_id*16+1], codeword_reg8[256*6+set_id*16+1], codeword_reg7[256*6+set_id*16+1], codeword_reg6[256*6+set_id*16+1], codeword_reg5[256*6+set_id*16+1], codeword_reg4[256*6+set_id*16+1], codeword_reg3[256*6+set_id*16+1], codeword_reg2[256*6+set_id*16+1], codeword_reg1[256*6+set_id*16+1], codeword_reg16[256*5+set_id*16+1], codeword_reg15[256*5+set_id*16+1], codeword_reg14[256*5+set_id*16+1], codeword_reg13[256*5+set_id*16+1], codeword_reg12[256*5+set_id*16+1], codeword_reg11[256*5+set_id*16+1], codeword_reg10[256*5+set_id*16+1], codeword_reg9[256*5+set_id*16+1], codeword_reg8[256*5+set_id*16+1], codeword_reg7[256*5+set_id*16+1], codeword_reg6[256*5+set_id*16+1], codeword_reg5[256*5+set_id*16+1], codeword_reg4[256*5+set_id*16+1], codeword_reg3[256*5+set_id*16+1], codeword_reg2[256*5+set_id*16+1], codeword_reg1[256*5+set_id*16+1], codeword_reg16[256*4+set_id*16+1], codeword_reg15[256*4+set_id*16+1], codeword_reg14[256*4+set_id*16+1], codeword_reg13[256*4+set_id*16+1], codeword_reg12[256*4+set_id*16+1], codeword_reg11[256*4+set_id*16+1], codeword_reg10[256*4+set_id*16+1], codeword_reg9[256*4+set_id*16+1], codeword_reg8[256*4+set_id*16+1], codeword_reg7[256*4+set_id*16+1], codeword_reg6[256*4+set_id*16+1], codeword_reg5[256*4+set_id*16+1], codeword_reg4[256*4+set_id*16+1], codeword_reg3[256*4+set_id*16+1], codeword_reg2[256*4+set_id*16+1], codeword_reg1[256*4+set_id*16+1], codeword_reg16[256*3+set_id*16+1], codeword_reg15[256*3+set_id*16+1], codeword_reg14[256*3+set_id*16+1], codeword_reg13[256*3+set_id*16+1], codeword_reg12[256*3+set_id*16+1], codeword_reg11[256*3+set_id*16+1], codeword_reg10[256*3+set_id*16+1], codeword_reg9[256*3+set_id*16+1], codeword_reg8[256*3+set_id*16+1], codeword_reg7[256*3+set_id*16+1], codeword_reg6[256*3+set_id*16+1], codeword_reg5[256*3+set_id*16+1], codeword_reg4[256*3+set_id*16+1], codeword_reg3[256*3+set_id*16+1], codeword_reg2[256*3+set_id*16+1], codeword_reg1[256*3+set_id*16+1], codeword_reg16[256*2+set_id*16+1], codeword_reg15[256*2+set_id*16+1], codeword_reg14[256*2+set_id*16+1], codeword_reg13[256*2+set_id*16+1], codeword_reg12[256*2+set_id*16+1], codeword_reg11[256*2+set_id*16+1], codeword_reg10[256*2+set_id*16+1], codeword_reg9[256*2+set_id*16+1], codeword_reg8[256*2+set_id*16+1], codeword_reg7[256*2+set_id*16+1], codeword_reg6[256*2+set_id*16+1], codeword_reg5[256*2+set_id*16+1], codeword_reg4[256*2+set_id*16+1], codeword_reg3[256*2+set_id*16+1], codeword_reg2[256*2+set_id*16+1], codeword_reg1[256*2+set_id*16+1], codeword_reg16[256*1+set_id*16+1], codeword_reg15[256*1+set_id*16+1], codeword_reg14[256*1+set_id*16+1], codeword_reg13[256*1+set_id*16+1], codeword_reg12[256*1+set_id*16+1], codeword_reg11[256*1+set_id*16+1], codeword_reg10[256*1+set_id*16+1], codeword_reg9[256*1+set_id*16+1], codeword_reg8[256*1+set_id*16+1], codeword_reg7[256*1+set_id*16+1], codeword_reg6[256*1+set_id*16+1], codeword_reg5[256*1+set_id*16+1], codeword_reg4[256*1+set_id*16+1], codeword_reg3[256*1+set_id*16+1], codeword_reg2[256*1+set_id*16+1], codeword_reg1[256*1+set_id*16+1], codeword_reg16[256*0+set_id*16+1], codeword_reg15[256*0+set_id*16+1], codeword_reg14[256*0+set_id*16+1], codeword_reg13[256*0+set_id*16+1], codeword_reg12[256*0+set_id*16+1], codeword_reg11[256*0+set_id*16+1], codeword_reg10[256*0+set_id*16+1], codeword_reg9[256*0+set_id*16+1], codeword_reg8[256*0+set_id*16+1], codeword_reg7[256*0+set_id*16+1], codeword_reg6[256*0+set_id*16+1], codeword_reg5[256*0+set_id*16+1], codeword_reg4[256*0+set_id*16+1], codeword_reg3[256*0+set_id*16+1], codeword_reg2[256*0+set_id*16+1], codeword_reg1[256*0+set_id*16+1]};
                            in_bits3  <= {codeword_reg16[256*14+set_id*16+2], codeword_reg15[256*14+set_id*16+2], codeword_reg14[256*14+set_id*16+2], codeword_reg13[256*14+set_id*16+2], codeword_reg12[256*14+set_id*16+2], codeword_reg11[256*14+set_id*16+2], codeword_reg10[256*14+set_id*16+2], codeword_reg9[256*14+set_id*16+2], codeword_reg8[256*14+set_id*16+2], codeword_reg7[256*14+set_id*16+2], codeword_reg6[256*14+set_id*16+2], codeword_reg5[256*14+set_id*16+2], codeword_reg4[256*14+set_id*16+2], codeword_reg3[256*14+set_id*16+2], codeword_reg2[256*14+set_id*16+2], codeword_reg1[256*14+set_id*16+2], codeword_reg16[256*13+set_id*16+2], codeword_reg15[256*13+set_id*16+2], codeword_reg14[256*13+set_id*16+2], codeword_reg13[256*13+set_id*16+2], codeword_reg12[256*13+set_id*16+2], codeword_reg11[256*13+set_id*16+2], codeword_reg10[256*13+set_id*16+2], codeword_reg9[256*13+set_id*16+2], codeword_reg8[256*13+set_id*16+2], codeword_reg7[256*13+set_id*16+2], codeword_reg6[256*13+set_id*16+2], codeword_reg5[256*13+set_id*16+2], codeword_reg4[256*13+set_id*16+2], codeword_reg3[256*13+set_id*16+2], codeword_reg2[256*13+set_id*16+2], codeword_reg1[256*13+set_id*16+2], codeword_reg16[256*12+set_id*16+2], codeword_reg15[256*12+set_id*16+2], codeword_reg14[256*12+set_id*16+2], codeword_reg13[256*12+set_id*16+2], codeword_reg12[256*12+set_id*16+2], codeword_reg11[256*12+set_id*16+2], codeword_reg10[256*12+set_id*16+2], codeword_reg9[256*12+set_id*16+2], codeword_reg8[256*12+set_id*16+2], codeword_reg7[256*12+set_id*16+2], codeword_reg6[256*12+set_id*16+2], codeword_reg5[256*12+set_id*16+2], codeword_reg4[256*12+set_id*16+2], codeword_reg3[256*12+set_id*16+2], codeword_reg2[256*12+set_id*16+2], codeword_reg1[256*12+set_id*16+2], codeword_reg16[256*11+set_id*16+2], codeword_reg15[256*11+set_id*16+2], codeword_reg14[256*11+set_id*16+2], codeword_reg13[256*11+set_id*16+2], codeword_reg12[256*11+set_id*16+2], codeword_reg11[256*11+set_id*16+2], codeword_reg10[256*11+set_id*16+2], codeword_reg9[256*11+set_id*16+2], codeword_reg8[256*11+set_id*16+2], codeword_reg7[256*11+set_id*16+2], codeword_reg6[256*11+set_id*16+2], codeword_reg5[256*11+set_id*16+2], codeword_reg4[256*11+set_id*16+2], codeword_reg3[256*11+set_id*16+2], codeword_reg2[256*11+set_id*16+2], codeword_reg1[256*11+set_id*16+2], codeword_reg16[256*10+set_id*16+2], codeword_reg15[256*10+set_id*16+2], codeword_reg14[256*10+set_id*16+2], codeword_reg13[256*10+set_id*16+2], codeword_reg12[256*10+set_id*16+2], codeword_reg11[256*10+set_id*16+2], codeword_reg10[256*10+set_id*16+2], codeword_reg9[256*10+set_id*16+2], codeword_reg8[256*10+set_id*16+2], codeword_reg7[256*10+set_id*16+2], codeword_reg6[256*10+set_id*16+2], codeword_reg5[256*10+set_id*16+2], codeword_reg4[256*10+set_id*16+2], codeword_reg3[256*10+set_id*16+2], codeword_reg2[256*10+set_id*16+2], codeword_reg1[256*10+set_id*16+2], codeword_reg16[256*9+set_id*16+2], codeword_reg15[256*9+set_id*16+2], codeword_reg14[256*9+set_id*16+2], codeword_reg13[256*9+set_id*16+2], codeword_reg12[256*9+set_id*16+2], codeword_reg11[256*9+set_id*16+2], codeword_reg10[256*9+set_id*16+2], codeword_reg9[256*9+set_id*16+2], codeword_reg8[256*9+set_id*16+2], codeword_reg7[256*9+set_id*16+2], codeword_reg6[256*9+set_id*16+2], codeword_reg5[256*9+set_id*16+2], codeword_reg4[256*9+set_id*16+2], codeword_reg3[256*9+set_id*16+2], codeword_reg2[256*9+set_id*16+2], codeword_reg1[256*9+set_id*16+2], codeword_reg16[256*8+set_id*16+2], codeword_reg15[256*8+set_id*16+2], codeword_reg14[256*8+set_id*16+2], codeword_reg13[256*8+set_id*16+2], codeword_reg12[256*8+set_id*16+2], codeword_reg11[256*8+set_id*16+2], codeword_reg10[256*8+set_id*16+2], codeword_reg9[256*8+set_id*16+2], codeword_reg8[256*8+set_id*16+2], codeword_reg7[256*8+set_id*16+2], codeword_reg6[256*8+set_id*16+2], codeword_reg5[256*8+set_id*16+2], codeword_reg4[256*8+set_id*16+2], codeword_reg3[256*8+set_id*16+2], codeword_reg2[256*8+set_id*16+2], codeword_reg1[256*8+set_id*16+2], codeword_reg16[256*7+set_id*16+2], codeword_reg15[256*7+set_id*16+2], codeword_reg14[256*7+set_id*16+2], codeword_reg13[256*7+set_id*16+2], codeword_reg12[256*7+set_id*16+2], codeword_reg11[256*7+set_id*16+2], codeword_reg10[256*7+set_id*16+2], codeword_reg9[256*7+set_id*16+2], codeword_reg8[256*7+set_id*16+2], codeword_reg7[256*7+set_id*16+2], codeword_reg6[256*7+set_id*16+2], codeword_reg5[256*7+set_id*16+2], codeword_reg4[256*7+set_id*16+2], codeword_reg3[256*7+set_id*16+2], codeword_reg2[256*7+set_id*16+2], codeword_reg1[256*7+set_id*16+2], codeword_reg16[256*6+set_id*16+2], codeword_reg15[256*6+set_id*16+2], codeword_reg14[256*6+set_id*16+2], codeword_reg13[256*6+set_id*16+2], codeword_reg12[256*6+set_id*16+2], codeword_reg11[256*6+set_id*16+2], codeword_reg10[256*6+set_id*16+2], codeword_reg9[256*6+set_id*16+2], codeword_reg8[256*6+set_id*16+2], codeword_reg7[256*6+set_id*16+2], codeword_reg6[256*6+set_id*16+2], codeword_reg5[256*6+set_id*16+2], codeword_reg4[256*6+set_id*16+2], codeword_reg3[256*6+set_id*16+2], codeword_reg2[256*6+set_id*16+2], codeword_reg1[256*6+set_id*16+2], codeword_reg16[256*5+set_id*16+2], codeword_reg15[256*5+set_id*16+2], codeword_reg14[256*5+set_id*16+2], codeword_reg13[256*5+set_id*16+2], codeword_reg12[256*5+set_id*16+2], codeword_reg11[256*5+set_id*16+2], codeword_reg10[256*5+set_id*16+2], codeword_reg9[256*5+set_id*16+2], codeword_reg8[256*5+set_id*16+2], codeword_reg7[256*5+set_id*16+2], codeword_reg6[256*5+set_id*16+2], codeword_reg5[256*5+set_id*16+2], codeword_reg4[256*5+set_id*16+2], codeword_reg3[256*5+set_id*16+2], codeword_reg2[256*5+set_id*16+2], codeword_reg1[256*5+set_id*16+2], codeword_reg16[256*4+set_id*16+2], codeword_reg15[256*4+set_id*16+2], codeword_reg14[256*4+set_id*16+2], codeword_reg13[256*4+set_id*16+2], codeword_reg12[256*4+set_id*16+2], codeword_reg11[256*4+set_id*16+2], codeword_reg10[256*4+set_id*16+2], codeword_reg9[256*4+set_id*16+2], codeword_reg8[256*4+set_id*16+2], codeword_reg7[256*4+set_id*16+2], codeword_reg6[256*4+set_id*16+2], codeword_reg5[256*4+set_id*16+2], codeword_reg4[256*4+set_id*16+2], codeword_reg3[256*4+set_id*16+2], codeword_reg2[256*4+set_id*16+2], codeword_reg1[256*4+set_id*16+2], codeword_reg16[256*3+set_id*16+2], codeword_reg15[256*3+set_id*16+2], codeword_reg14[256*3+set_id*16+2], codeword_reg13[256*3+set_id*16+2], codeword_reg12[256*3+set_id*16+2], codeword_reg11[256*3+set_id*16+2], codeword_reg10[256*3+set_id*16+2], codeword_reg9[256*3+set_id*16+2], codeword_reg8[256*3+set_id*16+2], codeword_reg7[256*3+set_id*16+2], codeword_reg6[256*3+set_id*16+2], codeword_reg5[256*3+set_id*16+2], codeword_reg4[256*3+set_id*16+2], codeword_reg3[256*3+set_id*16+2], codeword_reg2[256*3+set_id*16+2], codeword_reg1[256*3+set_id*16+2], codeword_reg16[256*2+set_id*16+2], codeword_reg15[256*2+set_id*16+2], codeword_reg14[256*2+set_id*16+2], codeword_reg13[256*2+set_id*16+2], codeword_reg12[256*2+set_id*16+2], codeword_reg11[256*2+set_id*16+2], codeword_reg10[256*2+set_id*16+2], codeword_reg9[256*2+set_id*16+2], codeword_reg8[256*2+set_id*16+2], codeword_reg7[256*2+set_id*16+2], codeword_reg6[256*2+set_id*16+2], codeword_reg5[256*2+set_id*16+2], codeword_reg4[256*2+set_id*16+2], codeword_reg3[256*2+set_id*16+2], codeword_reg2[256*2+set_id*16+2], codeword_reg1[256*2+set_id*16+2], codeword_reg16[256*1+set_id*16+2], codeword_reg15[256*1+set_id*16+2], codeword_reg14[256*1+set_id*16+2], codeword_reg13[256*1+set_id*16+2], codeword_reg12[256*1+set_id*16+2], codeword_reg11[256*1+set_id*16+2], codeword_reg10[256*1+set_id*16+2], codeword_reg9[256*1+set_id*16+2], codeword_reg8[256*1+set_id*16+2], codeword_reg7[256*1+set_id*16+2], codeword_reg6[256*1+set_id*16+2], codeword_reg5[256*1+set_id*16+2], codeword_reg4[256*1+set_id*16+2], codeword_reg3[256*1+set_id*16+2], codeword_reg2[256*1+set_id*16+2], codeword_reg1[256*1+set_id*16+2], codeword_reg16[256*0+set_id*16+2], codeword_reg15[256*0+set_id*16+2], codeword_reg14[256*0+set_id*16+2], codeword_reg13[256*0+set_id*16+2], codeword_reg12[256*0+set_id*16+2], codeword_reg11[256*0+set_id*16+2], codeword_reg10[256*0+set_id*16+2], codeword_reg9[256*0+set_id*16+2], codeword_reg8[256*0+set_id*16+2], codeword_reg7[256*0+set_id*16+2], codeword_reg6[256*0+set_id*16+2], codeword_reg5[256*0+set_id*16+2], codeword_reg4[256*0+set_id*16+2], codeword_reg3[256*0+set_id*16+2], codeword_reg2[256*0+set_id*16+2], codeword_reg1[256*0+set_id*16+2]};
                            in_bits4  <= {codeword_reg16[256*14+set_id*16+3], codeword_reg15[256*14+set_id*16+3], codeword_reg14[256*14+set_id*16+3], codeword_reg13[256*14+set_id*16+3], codeword_reg12[256*14+set_id*16+3], codeword_reg11[256*14+set_id*16+3], codeword_reg10[256*14+set_id*16+3], codeword_reg9[256*14+set_id*16+3], codeword_reg8[256*14+set_id*16+3], codeword_reg7[256*14+set_id*16+3], codeword_reg6[256*14+set_id*16+3], codeword_reg5[256*14+set_id*16+3], codeword_reg4[256*14+set_id*16+3], codeword_reg3[256*14+set_id*16+3], codeword_reg2[256*14+set_id*16+3], codeword_reg1[256*14+set_id*16+3], codeword_reg16[256*13+set_id*16+3], codeword_reg15[256*13+set_id*16+3], codeword_reg14[256*13+set_id*16+3], codeword_reg13[256*13+set_id*16+3], codeword_reg12[256*13+set_id*16+3], codeword_reg11[256*13+set_id*16+3], codeword_reg10[256*13+set_id*16+3], codeword_reg9[256*13+set_id*16+3], codeword_reg8[256*13+set_id*16+3], codeword_reg7[256*13+set_id*16+3], codeword_reg6[256*13+set_id*16+3], codeword_reg5[256*13+set_id*16+3], codeword_reg4[256*13+set_id*16+3], codeword_reg3[256*13+set_id*16+3], codeword_reg2[256*13+set_id*16+3], codeword_reg1[256*13+set_id*16+3], codeword_reg16[256*12+set_id*16+3], codeword_reg15[256*12+set_id*16+3], codeword_reg14[256*12+set_id*16+3], codeword_reg13[256*12+set_id*16+3], codeword_reg12[256*12+set_id*16+3], codeword_reg11[256*12+set_id*16+3], codeword_reg10[256*12+set_id*16+3], codeword_reg9[256*12+set_id*16+3], codeword_reg8[256*12+set_id*16+3], codeword_reg7[256*12+set_id*16+3], codeword_reg6[256*12+set_id*16+3], codeword_reg5[256*12+set_id*16+3], codeword_reg4[256*12+set_id*16+3], codeword_reg3[256*12+set_id*16+3], codeword_reg2[256*12+set_id*16+3], codeword_reg1[256*12+set_id*16+3], codeword_reg16[256*11+set_id*16+3], codeword_reg15[256*11+set_id*16+3], codeword_reg14[256*11+set_id*16+3], codeword_reg13[256*11+set_id*16+3], codeword_reg12[256*11+set_id*16+3], codeword_reg11[256*11+set_id*16+3], codeword_reg10[256*11+set_id*16+3], codeword_reg9[256*11+set_id*16+3], codeword_reg8[256*11+set_id*16+3], codeword_reg7[256*11+set_id*16+3], codeword_reg6[256*11+set_id*16+3], codeword_reg5[256*11+set_id*16+3], codeword_reg4[256*11+set_id*16+3], codeword_reg3[256*11+set_id*16+3], codeword_reg2[256*11+set_id*16+3], codeword_reg1[256*11+set_id*16+3], codeword_reg16[256*10+set_id*16+3], codeword_reg15[256*10+set_id*16+3], codeword_reg14[256*10+set_id*16+3], codeword_reg13[256*10+set_id*16+3], codeword_reg12[256*10+set_id*16+3], codeword_reg11[256*10+set_id*16+3], codeword_reg10[256*10+set_id*16+3], codeword_reg9[256*10+set_id*16+3], codeword_reg8[256*10+set_id*16+3], codeword_reg7[256*10+set_id*16+3], codeword_reg6[256*10+set_id*16+3], codeword_reg5[256*10+set_id*16+3], codeword_reg4[256*10+set_id*16+3], codeword_reg3[256*10+set_id*16+3], codeword_reg2[256*10+set_id*16+3], codeword_reg1[256*10+set_id*16+3], codeword_reg16[256*9+set_id*16+3], codeword_reg15[256*9+set_id*16+3], codeword_reg14[256*9+set_id*16+3], codeword_reg13[256*9+set_id*16+3], codeword_reg12[256*9+set_id*16+3], codeword_reg11[256*9+set_id*16+3], codeword_reg10[256*9+set_id*16+3], codeword_reg9[256*9+set_id*16+3], codeword_reg8[256*9+set_id*16+3], codeword_reg7[256*9+set_id*16+3], codeword_reg6[256*9+set_id*16+3], codeword_reg5[256*9+set_id*16+3], codeword_reg4[256*9+set_id*16+3], codeword_reg3[256*9+set_id*16+3], codeword_reg2[256*9+set_id*16+3], codeword_reg1[256*9+set_id*16+3], codeword_reg16[256*8+set_id*16+3], codeword_reg15[256*8+set_id*16+3], codeword_reg14[256*8+set_id*16+3], codeword_reg13[256*8+set_id*16+3], codeword_reg12[256*8+set_id*16+3], codeword_reg11[256*8+set_id*16+3], codeword_reg10[256*8+set_id*16+3], codeword_reg9[256*8+set_id*16+3], codeword_reg8[256*8+set_id*16+3], codeword_reg7[256*8+set_id*16+3], codeword_reg6[256*8+set_id*16+3], codeword_reg5[256*8+set_id*16+3], codeword_reg4[256*8+set_id*16+3], codeword_reg3[256*8+set_id*16+3], codeword_reg2[256*8+set_id*16+3], codeword_reg1[256*8+set_id*16+3], codeword_reg16[256*7+set_id*16+3], codeword_reg15[256*7+set_id*16+3], codeword_reg14[256*7+set_id*16+3], codeword_reg13[256*7+set_id*16+3], codeword_reg12[256*7+set_id*16+3], codeword_reg11[256*7+set_id*16+3], codeword_reg10[256*7+set_id*16+3], codeword_reg9[256*7+set_id*16+3], codeword_reg8[256*7+set_id*16+3], codeword_reg7[256*7+set_id*16+3], codeword_reg6[256*7+set_id*16+3], codeword_reg5[256*7+set_id*16+3], codeword_reg4[256*7+set_id*16+3], codeword_reg3[256*7+set_id*16+3], codeword_reg2[256*7+set_id*16+3], codeword_reg1[256*7+set_id*16+3], codeword_reg16[256*6+set_id*16+3], codeword_reg15[256*6+set_id*16+3], codeword_reg14[256*6+set_id*16+3], codeword_reg13[256*6+set_id*16+3], codeword_reg12[256*6+set_id*16+3], codeword_reg11[256*6+set_id*16+3], codeword_reg10[256*6+set_id*16+3], codeword_reg9[256*6+set_id*16+3], codeword_reg8[256*6+set_id*16+3], codeword_reg7[256*6+set_id*16+3], codeword_reg6[256*6+set_id*16+3], codeword_reg5[256*6+set_id*16+3], codeword_reg4[256*6+set_id*16+3], codeword_reg3[256*6+set_id*16+3], codeword_reg2[256*6+set_id*16+3], codeword_reg1[256*6+set_id*16+3], codeword_reg16[256*5+set_id*16+3], codeword_reg15[256*5+set_id*16+3], codeword_reg14[256*5+set_id*16+3], codeword_reg13[256*5+set_id*16+3], codeword_reg12[256*5+set_id*16+3], codeword_reg11[256*5+set_id*16+3], codeword_reg10[256*5+set_id*16+3], codeword_reg9[256*5+set_id*16+3], codeword_reg8[256*5+set_id*16+3], codeword_reg7[256*5+set_id*16+3], codeword_reg6[256*5+set_id*16+3], codeword_reg5[256*5+set_id*16+3], codeword_reg4[256*5+set_id*16+3], codeword_reg3[256*5+set_id*16+3], codeword_reg2[256*5+set_id*16+3], codeword_reg1[256*5+set_id*16+3], codeword_reg16[256*4+set_id*16+3], codeword_reg15[256*4+set_id*16+3], codeword_reg14[256*4+set_id*16+3], codeword_reg13[256*4+set_id*16+3], codeword_reg12[256*4+set_id*16+3], codeword_reg11[256*4+set_id*16+3], codeword_reg10[256*4+set_id*16+3], codeword_reg9[256*4+set_id*16+3], codeword_reg8[256*4+set_id*16+3], codeword_reg7[256*4+set_id*16+3], codeword_reg6[256*4+set_id*16+3], codeword_reg5[256*4+set_id*16+3], codeword_reg4[256*4+set_id*16+3], codeword_reg3[256*4+set_id*16+3], codeword_reg2[256*4+set_id*16+3], codeword_reg1[256*4+set_id*16+3], codeword_reg16[256*3+set_id*16+3], codeword_reg15[256*3+set_id*16+3], codeword_reg14[256*3+set_id*16+3], codeword_reg13[256*3+set_id*16+3], codeword_reg12[256*3+set_id*16+3], codeword_reg11[256*3+set_id*16+3], codeword_reg10[256*3+set_id*16+3], codeword_reg9[256*3+set_id*16+3], codeword_reg8[256*3+set_id*16+3], codeword_reg7[256*3+set_id*16+3], codeword_reg6[256*3+set_id*16+3], codeword_reg5[256*3+set_id*16+3], codeword_reg4[256*3+set_id*16+3], codeword_reg3[256*3+set_id*16+3], codeword_reg2[256*3+set_id*16+3], codeword_reg1[256*3+set_id*16+3], codeword_reg16[256*2+set_id*16+3], codeword_reg15[256*2+set_id*16+3], codeword_reg14[256*2+set_id*16+3], codeword_reg13[256*2+set_id*16+3], codeword_reg12[256*2+set_id*16+3], codeword_reg11[256*2+set_id*16+3], codeword_reg10[256*2+set_id*16+3], codeword_reg9[256*2+set_id*16+3], codeword_reg8[256*2+set_id*16+3], codeword_reg7[256*2+set_id*16+3], codeword_reg6[256*2+set_id*16+3], codeword_reg5[256*2+set_id*16+3], codeword_reg4[256*2+set_id*16+3], codeword_reg3[256*2+set_id*16+3], codeword_reg2[256*2+set_id*16+3], codeword_reg1[256*2+set_id*16+3], codeword_reg16[256*1+set_id*16+3], codeword_reg15[256*1+set_id*16+3], codeword_reg14[256*1+set_id*16+3], codeword_reg13[256*1+set_id*16+3], codeword_reg12[256*1+set_id*16+3], codeword_reg11[256*1+set_id*16+3], codeword_reg10[256*1+set_id*16+3], codeword_reg9[256*1+set_id*16+3], codeword_reg8[256*1+set_id*16+3], codeword_reg7[256*1+set_id*16+3], codeword_reg6[256*1+set_id*16+3], codeword_reg5[256*1+set_id*16+3], codeword_reg4[256*1+set_id*16+3], codeword_reg3[256*1+set_id*16+3], codeword_reg2[256*1+set_id*16+3], codeword_reg1[256*1+set_id*16+3], codeword_reg16[256*0+set_id*16+3], codeword_reg15[256*0+set_id*16+3], codeword_reg14[256*0+set_id*16+3], codeword_reg13[256*0+set_id*16+3], codeword_reg12[256*0+set_id*16+3], codeword_reg11[256*0+set_id*16+3], codeword_reg10[256*0+set_id*16+3], codeword_reg9[256*0+set_id*16+3], codeword_reg8[256*0+set_id*16+3], codeword_reg7[256*0+set_id*16+3], codeword_reg6[256*0+set_id*16+3], codeword_reg5[256*0+set_id*16+3], codeword_reg4[256*0+set_id*16+3], codeword_reg3[256*0+set_id*16+3], codeword_reg2[256*0+set_id*16+3], codeword_reg1[256*0+set_id*16+3]};
                            in_bits5  <= {codeword_reg16[256*14+set_id*16+4], codeword_reg15[256*14+set_id*16+4], codeword_reg14[256*14+set_id*16+4], codeword_reg13[256*14+set_id*16+4], codeword_reg12[256*14+set_id*16+4], codeword_reg11[256*14+set_id*16+4], codeword_reg10[256*14+set_id*16+4], codeword_reg9[256*14+set_id*16+4], codeword_reg8[256*14+set_id*16+4], codeword_reg7[256*14+set_id*16+4], codeword_reg6[256*14+set_id*16+4], codeword_reg5[256*14+set_id*16+4], codeword_reg4[256*14+set_id*16+4], codeword_reg3[256*14+set_id*16+4], codeword_reg2[256*14+set_id*16+4], codeword_reg1[256*14+set_id*16+4], codeword_reg16[256*13+set_id*16+4], codeword_reg15[256*13+set_id*16+4], codeword_reg14[256*13+set_id*16+4], codeword_reg13[256*13+set_id*16+4], codeword_reg12[256*13+set_id*16+4], codeword_reg11[256*13+set_id*16+4], codeword_reg10[256*13+set_id*16+4], codeword_reg9[256*13+set_id*16+4], codeword_reg8[256*13+set_id*16+4], codeword_reg7[256*13+set_id*16+4], codeword_reg6[256*13+set_id*16+4], codeword_reg5[256*13+set_id*16+4], codeword_reg4[256*13+set_id*16+4], codeword_reg3[256*13+set_id*16+4], codeword_reg2[256*13+set_id*16+4], codeword_reg1[256*13+set_id*16+4], codeword_reg16[256*12+set_id*16+4], codeword_reg15[256*12+set_id*16+4], codeword_reg14[256*12+set_id*16+4], codeword_reg13[256*12+set_id*16+4], codeword_reg12[256*12+set_id*16+4], codeword_reg11[256*12+set_id*16+4], codeword_reg10[256*12+set_id*16+4], codeword_reg9[256*12+set_id*16+4], codeword_reg8[256*12+set_id*16+4], codeword_reg7[256*12+set_id*16+4], codeword_reg6[256*12+set_id*16+4], codeword_reg5[256*12+set_id*16+4], codeword_reg4[256*12+set_id*16+4], codeword_reg3[256*12+set_id*16+4], codeword_reg2[256*12+set_id*16+4], codeword_reg1[256*12+set_id*16+4], codeword_reg16[256*11+set_id*16+4], codeword_reg15[256*11+set_id*16+4], codeword_reg14[256*11+set_id*16+4], codeword_reg13[256*11+set_id*16+4], codeword_reg12[256*11+set_id*16+4], codeword_reg11[256*11+set_id*16+4], codeword_reg10[256*11+set_id*16+4], codeword_reg9[256*11+set_id*16+4], codeword_reg8[256*11+set_id*16+4], codeword_reg7[256*11+set_id*16+4], codeword_reg6[256*11+set_id*16+4], codeword_reg5[256*11+set_id*16+4], codeword_reg4[256*11+set_id*16+4], codeword_reg3[256*11+set_id*16+4], codeword_reg2[256*11+set_id*16+4], codeword_reg1[256*11+set_id*16+4], codeword_reg16[256*10+set_id*16+4], codeword_reg15[256*10+set_id*16+4], codeword_reg14[256*10+set_id*16+4], codeword_reg13[256*10+set_id*16+4], codeword_reg12[256*10+set_id*16+4], codeword_reg11[256*10+set_id*16+4], codeword_reg10[256*10+set_id*16+4], codeword_reg9[256*10+set_id*16+4], codeword_reg8[256*10+set_id*16+4], codeword_reg7[256*10+set_id*16+4], codeword_reg6[256*10+set_id*16+4], codeword_reg5[256*10+set_id*16+4], codeword_reg4[256*10+set_id*16+4], codeword_reg3[256*10+set_id*16+4], codeword_reg2[256*10+set_id*16+4], codeword_reg1[256*10+set_id*16+4], codeword_reg16[256*9+set_id*16+4], codeword_reg15[256*9+set_id*16+4], codeword_reg14[256*9+set_id*16+4], codeword_reg13[256*9+set_id*16+4], codeword_reg12[256*9+set_id*16+4], codeword_reg11[256*9+set_id*16+4], codeword_reg10[256*9+set_id*16+4], codeword_reg9[256*9+set_id*16+4], codeword_reg8[256*9+set_id*16+4], codeword_reg7[256*9+set_id*16+4], codeword_reg6[256*9+set_id*16+4], codeword_reg5[256*9+set_id*16+4], codeword_reg4[256*9+set_id*16+4], codeword_reg3[256*9+set_id*16+4], codeword_reg2[256*9+set_id*16+4], codeword_reg1[256*9+set_id*16+4], codeword_reg16[256*8+set_id*16+4], codeword_reg15[256*8+set_id*16+4], codeword_reg14[256*8+set_id*16+4], codeword_reg13[256*8+set_id*16+4], codeword_reg12[256*8+set_id*16+4], codeword_reg11[256*8+set_id*16+4], codeword_reg10[256*8+set_id*16+4], codeword_reg9[256*8+set_id*16+4], codeword_reg8[256*8+set_id*16+4], codeword_reg7[256*8+set_id*16+4], codeword_reg6[256*8+set_id*16+4], codeword_reg5[256*8+set_id*16+4], codeword_reg4[256*8+set_id*16+4], codeword_reg3[256*8+set_id*16+4], codeword_reg2[256*8+set_id*16+4], codeword_reg1[256*8+set_id*16+4], codeword_reg16[256*7+set_id*16+4], codeword_reg15[256*7+set_id*16+4], codeword_reg14[256*7+set_id*16+4], codeword_reg13[256*7+set_id*16+4], codeword_reg12[256*7+set_id*16+4], codeword_reg11[256*7+set_id*16+4], codeword_reg10[256*7+set_id*16+4], codeword_reg9[256*7+set_id*16+4], codeword_reg8[256*7+set_id*16+4], codeword_reg7[256*7+set_id*16+4], codeword_reg6[256*7+set_id*16+4], codeword_reg5[256*7+set_id*16+4], codeword_reg4[256*7+set_id*16+4], codeword_reg3[256*7+set_id*16+4], codeword_reg2[256*7+set_id*16+4], codeword_reg1[256*7+set_id*16+4], codeword_reg16[256*6+set_id*16+4], codeword_reg15[256*6+set_id*16+4], codeword_reg14[256*6+set_id*16+4], codeword_reg13[256*6+set_id*16+4], codeword_reg12[256*6+set_id*16+4], codeword_reg11[256*6+set_id*16+4], codeword_reg10[256*6+set_id*16+4], codeword_reg9[256*6+set_id*16+4], codeword_reg8[256*6+set_id*16+4], codeword_reg7[256*6+set_id*16+4], codeword_reg6[256*6+set_id*16+4], codeword_reg5[256*6+set_id*16+4], codeword_reg4[256*6+set_id*16+4], codeword_reg3[256*6+set_id*16+4], codeword_reg2[256*6+set_id*16+4], codeword_reg1[256*6+set_id*16+4], codeword_reg16[256*5+set_id*16+4], codeword_reg15[256*5+set_id*16+4], codeword_reg14[256*5+set_id*16+4], codeword_reg13[256*5+set_id*16+4], codeword_reg12[256*5+set_id*16+4], codeword_reg11[256*5+set_id*16+4], codeword_reg10[256*5+set_id*16+4], codeword_reg9[256*5+set_id*16+4], codeword_reg8[256*5+set_id*16+4], codeword_reg7[256*5+set_id*16+4], codeword_reg6[256*5+set_id*16+4], codeword_reg5[256*5+set_id*16+4], codeword_reg4[256*5+set_id*16+4], codeword_reg3[256*5+set_id*16+4], codeword_reg2[256*5+set_id*16+4], codeword_reg1[256*5+set_id*16+4], codeword_reg16[256*4+set_id*16+4], codeword_reg15[256*4+set_id*16+4], codeword_reg14[256*4+set_id*16+4], codeword_reg13[256*4+set_id*16+4], codeword_reg12[256*4+set_id*16+4], codeword_reg11[256*4+set_id*16+4], codeword_reg10[256*4+set_id*16+4], codeword_reg9[256*4+set_id*16+4], codeword_reg8[256*4+set_id*16+4], codeword_reg7[256*4+set_id*16+4], codeword_reg6[256*4+set_id*16+4], codeword_reg5[256*4+set_id*16+4], codeword_reg4[256*4+set_id*16+4], codeword_reg3[256*4+set_id*16+4], codeword_reg2[256*4+set_id*16+4], codeword_reg1[256*4+set_id*16+4], codeword_reg16[256*3+set_id*16+4], codeword_reg15[256*3+set_id*16+4], codeword_reg14[256*3+set_id*16+4], codeword_reg13[256*3+set_id*16+4], codeword_reg12[256*3+set_id*16+4], codeword_reg11[256*3+set_id*16+4], codeword_reg10[256*3+set_id*16+4], codeword_reg9[256*3+set_id*16+4], codeword_reg8[256*3+set_id*16+4], codeword_reg7[256*3+set_id*16+4], codeword_reg6[256*3+set_id*16+4], codeword_reg5[256*3+set_id*16+4], codeword_reg4[256*3+set_id*16+4], codeword_reg3[256*3+set_id*16+4], codeword_reg2[256*3+set_id*16+4], codeword_reg1[256*3+set_id*16+4], codeword_reg16[256*2+set_id*16+4], codeword_reg15[256*2+set_id*16+4], codeword_reg14[256*2+set_id*16+4], codeword_reg13[256*2+set_id*16+4], codeword_reg12[256*2+set_id*16+4], codeword_reg11[256*2+set_id*16+4], codeword_reg10[256*2+set_id*16+4], codeword_reg9[256*2+set_id*16+4], codeword_reg8[256*2+set_id*16+4], codeword_reg7[256*2+set_id*16+4], codeword_reg6[256*2+set_id*16+4], codeword_reg5[256*2+set_id*16+4], codeword_reg4[256*2+set_id*16+4], codeword_reg3[256*2+set_id*16+4], codeword_reg2[256*2+set_id*16+4], codeword_reg1[256*2+set_id*16+4], codeword_reg16[256*1+set_id*16+4], codeword_reg15[256*1+set_id*16+4], codeword_reg14[256*1+set_id*16+4], codeword_reg13[256*1+set_id*16+4], codeword_reg12[256*1+set_id*16+4], codeword_reg11[256*1+set_id*16+4], codeword_reg10[256*1+set_id*16+4], codeword_reg9[256*1+set_id*16+4], codeword_reg8[256*1+set_id*16+4], codeword_reg7[256*1+set_id*16+4], codeword_reg6[256*1+set_id*16+4], codeword_reg5[256*1+set_id*16+4], codeword_reg4[256*1+set_id*16+4], codeword_reg3[256*1+set_id*16+4], codeword_reg2[256*1+set_id*16+4], codeword_reg1[256*1+set_id*16+4], codeword_reg16[256*0+set_id*16+4], codeword_reg15[256*0+set_id*16+4], codeword_reg14[256*0+set_id*16+4], codeword_reg13[256*0+set_id*16+4], codeword_reg12[256*0+set_id*16+4], codeword_reg11[256*0+set_id*16+4], codeword_reg10[256*0+set_id*16+4], codeword_reg9[256*0+set_id*16+4], codeword_reg8[256*0+set_id*16+4], codeword_reg7[256*0+set_id*16+4], codeword_reg6[256*0+set_id*16+4], codeword_reg5[256*0+set_id*16+4], codeword_reg4[256*0+set_id*16+4], codeword_reg3[256*0+set_id*16+4], codeword_reg2[256*0+set_id*16+4], codeword_reg1[256*0+set_id*16+4]};
                            in_bits6  <= {codeword_reg16[256*14+set_id*16+5], codeword_reg15[256*14+set_id*16+5], codeword_reg14[256*14+set_id*16+5], codeword_reg13[256*14+set_id*16+5], codeword_reg12[256*14+set_id*16+5], codeword_reg11[256*14+set_id*16+5], codeword_reg10[256*14+set_id*16+5], codeword_reg9[256*14+set_id*16+5], codeword_reg8[256*14+set_id*16+5], codeword_reg7[256*14+set_id*16+5], codeword_reg6[256*14+set_id*16+5], codeword_reg5[256*14+set_id*16+5], codeword_reg4[256*14+set_id*16+5], codeword_reg3[256*14+set_id*16+5], codeword_reg2[256*14+set_id*16+5], codeword_reg1[256*14+set_id*16+5], codeword_reg16[256*13+set_id*16+5], codeword_reg15[256*13+set_id*16+5], codeword_reg14[256*13+set_id*16+5], codeword_reg13[256*13+set_id*16+5], codeword_reg12[256*13+set_id*16+5], codeword_reg11[256*13+set_id*16+5], codeword_reg10[256*13+set_id*16+5], codeword_reg9[256*13+set_id*16+5], codeword_reg8[256*13+set_id*16+5], codeword_reg7[256*13+set_id*16+5], codeword_reg6[256*13+set_id*16+5], codeword_reg5[256*13+set_id*16+5], codeword_reg4[256*13+set_id*16+5], codeword_reg3[256*13+set_id*16+5], codeword_reg2[256*13+set_id*16+5], codeword_reg1[256*13+set_id*16+5], codeword_reg16[256*12+set_id*16+5], codeword_reg15[256*12+set_id*16+5], codeword_reg14[256*12+set_id*16+5], codeword_reg13[256*12+set_id*16+5], codeword_reg12[256*12+set_id*16+5], codeword_reg11[256*12+set_id*16+5], codeword_reg10[256*12+set_id*16+5], codeword_reg9[256*12+set_id*16+5], codeword_reg8[256*12+set_id*16+5], codeword_reg7[256*12+set_id*16+5], codeword_reg6[256*12+set_id*16+5], codeword_reg5[256*12+set_id*16+5], codeword_reg4[256*12+set_id*16+5], codeword_reg3[256*12+set_id*16+5], codeword_reg2[256*12+set_id*16+5], codeword_reg1[256*12+set_id*16+5], codeword_reg16[256*11+set_id*16+5], codeword_reg15[256*11+set_id*16+5], codeword_reg14[256*11+set_id*16+5], codeword_reg13[256*11+set_id*16+5], codeword_reg12[256*11+set_id*16+5], codeword_reg11[256*11+set_id*16+5], codeword_reg10[256*11+set_id*16+5], codeword_reg9[256*11+set_id*16+5], codeword_reg8[256*11+set_id*16+5], codeword_reg7[256*11+set_id*16+5], codeword_reg6[256*11+set_id*16+5], codeword_reg5[256*11+set_id*16+5], codeword_reg4[256*11+set_id*16+5], codeword_reg3[256*11+set_id*16+5], codeword_reg2[256*11+set_id*16+5], codeword_reg1[256*11+set_id*16+5], codeword_reg16[256*10+set_id*16+5], codeword_reg15[256*10+set_id*16+5], codeword_reg14[256*10+set_id*16+5], codeword_reg13[256*10+set_id*16+5], codeword_reg12[256*10+set_id*16+5], codeword_reg11[256*10+set_id*16+5], codeword_reg10[256*10+set_id*16+5], codeword_reg9[256*10+set_id*16+5], codeword_reg8[256*10+set_id*16+5], codeword_reg7[256*10+set_id*16+5], codeword_reg6[256*10+set_id*16+5], codeword_reg5[256*10+set_id*16+5], codeword_reg4[256*10+set_id*16+5], codeword_reg3[256*10+set_id*16+5], codeword_reg2[256*10+set_id*16+5], codeword_reg1[256*10+set_id*16+5], codeword_reg16[256*9+set_id*16+5], codeword_reg15[256*9+set_id*16+5], codeword_reg14[256*9+set_id*16+5], codeword_reg13[256*9+set_id*16+5], codeword_reg12[256*9+set_id*16+5], codeword_reg11[256*9+set_id*16+5], codeword_reg10[256*9+set_id*16+5], codeword_reg9[256*9+set_id*16+5], codeword_reg8[256*9+set_id*16+5], codeword_reg7[256*9+set_id*16+5], codeword_reg6[256*9+set_id*16+5], codeword_reg5[256*9+set_id*16+5], codeword_reg4[256*9+set_id*16+5], codeword_reg3[256*9+set_id*16+5], codeword_reg2[256*9+set_id*16+5], codeword_reg1[256*9+set_id*16+5], codeword_reg16[256*8+set_id*16+5], codeword_reg15[256*8+set_id*16+5], codeword_reg14[256*8+set_id*16+5], codeword_reg13[256*8+set_id*16+5], codeword_reg12[256*8+set_id*16+5], codeword_reg11[256*8+set_id*16+5], codeword_reg10[256*8+set_id*16+5], codeword_reg9[256*8+set_id*16+5], codeword_reg8[256*8+set_id*16+5], codeword_reg7[256*8+set_id*16+5], codeword_reg6[256*8+set_id*16+5], codeword_reg5[256*8+set_id*16+5], codeword_reg4[256*8+set_id*16+5], codeword_reg3[256*8+set_id*16+5], codeword_reg2[256*8+set_id*16+5], codeword_reg1[256*8+set_id*16+5], codeword_reg16[256*7+set_id*16+5], codeword_reg15[256*7+set_id*16+5], codeword_reg14[256*7+set_id*16+5], codeword_reg13[256*7+set_id*16+5], codeword_reg12[256*7+set_id*16+5], codeword_reg11[256*7+set_id*16+5], codeword_reg10[256*7+set_id*16+5], codeword_reg9[256*7+set_id*16+5], codeword_reg8[256*7+set_id*16+5], codeword_reg7[256*7+set_id*16+5], codeword_reg6[256*7+set_id*16+5], codeword_reg5[256*7+set_id*16+5], codeword_reg4[256*7+set_id*16+5], codeword_reg3[256*7+set_id*16+5], codeword_reg2[256*7+set_id*16+5], codeword_reg1[256*7+set_id*16+5], codeword_reg16[256*6+set_id*16+5], codeword_reg15[256*6+set_id*16+5], codeword_reg14[256*6+set_id*16+5], codeword_reg13[256*6+set_id*16+5], codeword_reg12[256*6+set_id*16+5], codeword_reg11[256*6+set_id*16+5], codeword_reg10[256*6+set_id*16+5], codeword_reg9[256*6+set_id*16+5], codeword_reg8[256*6+set_id*16+5], codeword_reg7[256*6+set_id*16+5], codeword_reg6[256*6+set_id*16+5], codeword_reg5[256*6+set_id*16+5], codeword_reg4[256*6+set_id*16+5], codeword_reg3[256*6+set_id*16+5], codeword_reg2[256*6+set_id*16+5], codeword_reg1[256*6+set_id*16+5], codeword_reg16[256*5+set_id*16+5], codeword_reg15[256*5+set_id*16+5], codeword_reg14[256*5+set_id*16+5], codeword_reg13[256*5+set_id*16+5], codeword_reg12[256*5+set_id*16+5], codeword_reg11[256*5+set_id*16+5], codeword_reg10[256*5+set_id*16+5], codeword_reg9[256*5+set_id*16+5], codeword_reg8[256*5+set_id*16+5], codeword_reg7[256*5+set_id*16+5], codeword_reg6[256*5+set_id*16+5], codeword_reg5[256*5+set_id*16+5], codeword_reg4[256*5+set_id*16+5], codeword_reg3[256*5+set_id*16+5], codeword_reg2[256*5+set_id*16+5], codeword_reg1[256*5+set_id*16+5], codeword_reg16[256*4+set_id*16+5], codeword_reg15[256*4+set_id*16+5], codeword_reg14[256*4+set_id*16+5], codeword_reg13[256*4+set_id*16+5], codeword_reg12[256*4+set_id*16+5], codeword_reg11[256*4+set_id*16+5], codeword_reg10[256*4+set_id*16+5], codeword_reg9[256*4+set_id*16+5], codeword_reg8[256*4+set_id*16+5], codeword_reg7[256*4+set_id*16+5], codeword_reg6[256*4+set_id*16+5], codeword_reg5[256*4+set_id*16+5], codeword_reg4[256*4+set_id*16+5], codeword_reg3[256*4+set_id*16+5], codeword_reg2[256*4+set_id*16+5], codeword_reg1[256*4+set_id*16+5], codeword_reg16[256*3+set_id*16+5], codeword_reg15[256*3+set_id*16+5], codeword_reg14[256*3+set_id*16+5], codeword_reg13[256*3+set_id*16+5], codeword_reg12[256*3+set_id*16+5], codeword_reg11[256*3+set_id*16+5], codeword_reg10[256*3+set_id*16+5], codeword_reg9[256*3+set_id*16+5], codeword_reg8[256*3+set_id*16+5], codeword_reg7[256*3+set_id*16+5], codeword_reg6[256*3+set_id*16+5], codeword_reg5[256*3+set_id*16+5], codeword_reg4[256*3+set_id*16+5], codeword_reg3[256*3+set_id*16+5], codeword_reg2[256*3+set_id*16+5], codeword_reg1[256*3+set_id*16+5], codeword_reg16[256*2+set_id*16+5], codeword_reg15[256*2+set_id*16+5], codeword_reg14[256*2+set_id*16+5], codeword_reg13[256*2+set_id*16+5], codeword_reg12[256*2+set_id*16+5], codeword_reg11[256*2+set_id*16+5], codeword_reg10[256*2+set_id*16+5], codeword_reg9[256*2+set_id*16+5], codeword_reg8[256*2+set_id*16+5], codeword_reg7[256*2+set_id*16+5], codeword_reg6[256*2+set_id*16+5], codeword_reg5[256*2+set_id*16+5], codeword_reg4[256*2+set_id*16+5], codeword_reg3[256*2+set_id*16+5], codeword_reg2[256*2+set_id*16+5], codeword_reg1[256*2+set_id*16+5], codeword_reg16[256*1+set_id*16+5], codeword_reg15[256*1+set_id*16+5], codeword_reg14[256*1+set_id*16+5], codeword_reg13[256*1+set_id*16+5], codeword_reg12[256*1+set_id*16+5], codeword_reg11[256*1+set_id*16+5], codeword_reg10[256*1+set_id*16+5], codeword_reg9[256*1+set_id*16+5], codeword_reg8[256*1+set_id*16+5], codeword_reg7[256*1+set_id*16+5], codeword_reg6[256*1+set_id*16+5], codeword_reg5[256*1+set_id*16+5], codeword_reg4[256*1+set_id*16+5], codeword_reg3[256*1+set_id*16+5], codeword_reg2[256*1+set_id*16+5], codeword_reg1[256*1+set_id*16+5], codeword_reg16[256*0+set_id*16+5], codeword_reg15[256*0+set_id*16+5], codeword_reg14[256*0+set_id*16+5], codeword_reg13[256*0+set_id*16+5], codeword_reg12[256*0+set_id*16+5], codeword_reg11[256*0+set_id*16+5], codeword_reg10[256*0+set_id*16+5], codeword_reg9[256*0+set_id*16+5], codeword_reg8[256*0+set_id*16+5], codeword_reg7[256*0+set_id*16+5], codeword_reg6[256*0+set_id*16+5], codeword_reg5[256*0+set_id*16+5], codeword_reg4[256*0+set_id*16+5], codeword_reg3[256*0+set_id*16+5], codeword_reg2[256*0+set_id*16+5], codeword_reg1[256*0+set_id*16+5]};
                            in_bits7  <= {codeword_reg16[256*14+set_id*16+6], codeword_reg15[256*14+set_id*16+6], codeword_reg14[256*14+set_id*16+6], codeword_reg13[256*14+set_id*16+6], codeword_reg12[256*14+set_id*16+6], codeword_reg11[256*14+set_id*16+6], codeword_reg10[256*14+set_id*16+6], codeword_reg9[256*14+set_id*16+6], codeword_reg8[256*14+set_id*16+6], codeword_reg7[256*14+set_id*16+6], codeword_reg6[256*14+set_id*16+6], codeword_reg5[256*14+set_id*16+6], codeword_reg4[256*14+set_id*16+6], codeword_reg3[256*14+set_id*16+6], codeword_reg2[256*14+set_id*16+6], codeword_reg1[256*14+set_id*16+6], codeword_reg16[256*13+set_id*16+6], codeword_reg15[256*13+set_id*16+6], codeword_reg14[256*13+set_id*16+6], codeword_reg13[256*13+set_id*16+6], codeword_reg12[256*13+set_id*16+6], codeword_reg11[256*13+set_id*16+6], codeword_reg10[256*13+set_id*16+6], codeword_reg9[256*13+set_id*16+6], codeword_reg8[256*13+set_id*16+6], codeword_reg7[256*13+set_id*16+6], codeword_reg6[256*13+set_id*16+6], codeword_reg5[256*13+set_id*16+6], codeword_reg4[256*13+set_id*16+6], codeword_reg3[256*13+set_id*16+6], codeword_reg2[256*13+set_id*16+6], codeword_reg1[256*13+set_id*16+6], codeword_reg16[256*12+set_id*16+6], codeword_reg15[256*12+set_id*16+6], codeword_reg14[256*12+set_id*16+6], codeword_reg13[256*12+set_id*16+6], codeword_reg12[256*12+set_id*16+6], codeword_reg11[256*12+set_id*16+6], codeword_reg10[256*12+set_id*16+6], codeword_reg9[256*12+set_id*16+6], codeword_reg8[256*12+set_id*16+6], codeword_reg7[256*12+set_id*16+6], codeword_reg6[256*12+set_id*16+6], codeword_reg5[256*12+set_id*16+6], codeword_reg4[256*12+set_id*16+6], codeword_reg3[256*12+set_id*16+6], codeword_reg2[256*12+set_id*16+6], codeword_reg1[256*12+set_id*16+6], codeword_reg16[256*11+set_id*16+6], codeword_reg15[256*11+set_id*16+6], codeword_reg14[256*11+set_id*16+6], codeword_reg13[256*11+set_id*16+6], codeword_reg12[256*11+set_id*16+6], codeword_reg11[256*11+set_id*16+6], codeword_reg10[256*11+set_id*16+6], codeword_reg9[256*11+set_id*16+6], codeword_reg8[256*11+set_id*16+6], codeword_reg7[256*11+set_id*16+6], codeword_reg6[256*11+set_id*16+6], codeword_reg5[256*11+set_id*16+6], codeword_reg4[256*11+set_id*16+6], codeword_reg3[256*11+set_id*16+6], codeword_reg2[256*11+set_id*16+6], codeword_reg1[256*11+set_id*16+6], codeword_reg16[256*10+set_id*16+6], codeword_reg15[256*10+set_id*16+6], codeword_reg14[256*10+set_id*16+6], codeword_reg13[256*10+set_id*16+6], codeword_reg12[256*10+set_id*16+6], codeword_reg11[256*10+set_id*16+6], codeword_reg10[256*10+set_id*16+6], codeword_reg9[256*10+set_id*16+6], codeword_reg8[256*10+set_id*16+6], codeword_reg7[256*10+set_id*16+6], codeword_reg6[256*10+set_id*16+6], codeword_reg5[256*10+set_id*16+6], codeword_reg4[256*10+set_id*16+6], codeword_reg3[256*10+set_id*16+6], codeword_reg2[256*10+set_id*16+6], codeword_reg1[256*10+set_id*16+6], codeword_reg16[256*9+set_id*16+6], codeword_reg15[256*9+set_id*16+6], codeword_reg14[256*9+set_id*16+6], codeword_reg13[256*9+set_id*16+6], codeword_reg12[256*9+set_id*16+6], codeword_reg11[256*9+set_id*16+6], codeword_reg10[256*9+set_id*16+6], codeword_reg9[256*9+set_id*16+6], codeword_reg8[256*9+set_id*16+6], codeword_reg7[256*9+set_id*16+6], codeword_reg6[256*9+set_id*16+6], codeword_reg5[256*9+set_id*16+6], codeword_reg4[256*9+set_id*16+6], codeword_reg3[256*9+set_id*16+6], codeword_reg2[256*9+set_id*16+6], codeword_reg1[256*9+set_id*16+6], codeword_reg16[256*8+set_id*16+6], codeword_reg15[256*8+set_id*16+6], codeword_reg14[256*8+set_id*16+6], codeword_reg13[256*8+set_id*16+6], codeword_reg12[256*8+set_id*16+6], codeword_reg11[256*8+set_id*16+6], codeword_reg10[256*8+set_id*16+6], codeword_reg9[256*8+set_id*16+6], codeword_reg8[256*8+set_id*16+6], codeword_reg7[256*8+set_id*16+6], codeword_reg6[256*8+set_id*16+6], codeword_reg5[256*8+set_id*16+6], codeword_reg4[256*8+set_id*16+6], codeword_reg3[256*8+set_id*16+6], codeword_reg2[256*8+set_id*16+6], codeword_reg1[256*8+set_id*16+6], codeword_reg16[256*7+set_id*16+6], codeword_reg15[256*7+set_id*16+6], codeword_reg14[256*7+set_id*16+6], codeword_reg13[256*7+set_id*16+6], codeword_reg12[256*7+set_id*16+6], codeword_reg11[256*7+set_id*16+6], codeword_reg10[256*7+set_id*16+6], codeword_reg9[256*7+set_id*16+6], codeword_reg8[256*7+set_id*16+6], codeword_reg7[256*7+set_id*16+6], codeword_reg6[256*7+set_id*16+6], codeword_reg5[256*7+set_id*16+6], codeword_reg4[256*7+set_id*16+6], codeword_reg3[256*7+set_id*16+6], codeword_reg2[256*7+set_id*16+6], codeword_reg1[256*7+set_id*16+6], codeword_reg16[256*6+set_id*16+6], codeword_reg15[256*6+set_id*16+6], codeword_reg14[256*6+set_id*16+6], codeword_reg13[256*6+set_id*16+6], codeword_reg12[256*6+set_id*16+6], codeword_reg11[256*6+set_id*16+6], codeword_reg10[256*6+set_id*16+6], codeword_reg9[256*6+set_id*16+6], codeword_reg8[256*6+set_id*16+6], codeword_reg7[256*6+set_id*16+6], codeword_reg6[256*6+set_id*16+6], codeword_reg5[256*6+set_id*16+6], codeword_reg4[256*6+set_id*16+6], codeword_reg3[256*6+set_id*16+6], codeword_reg2[256*6+set_id*16+6], codeword_reg1[256*6+set_id*16+6], codeword_reg16[256*5+set_id*16+6], codeword_reg15[256*5+set_id*16+6], codeword_reg14[256*5+set_id*16+6], codeword_reg13[256*5+set_id*16+6], codeword_reg12[256*5+set_id*16+6], codeword_reg11[256*5+set_id*16+6], codeword_reg10[256*5+set_id*16+6], codeword_reg9[256*5+set_id*16+6], codeword_reg8[256*5+set_id*16+6], codeword_reg7[256*5+set_id*16+6], codeword_reg6[256*5+set_id*16+6], codeword_reg5[256*5+set_id*16+6], codeword_reg4[256*5+set_id*16+6], codeword_reg3[256*5+set_id*16+6], codeword_reg2[256*5+set_id*16+6], codeword_reg1[256*5+set_id*16+6], codeword_reg16[256*4+set_id*16+6], codeword_reg15[256*4+set_id*16+6], codeword_reg14[256*4+set_id*16+6], codeword_reg13[256*4+set_id*16+6], codeword_reg12[256*4+set_id*16+6], codeword_reg11[256*4+set_id*16+6], codeword_reg10[256*4+set_id*16+6], codeword_reg9[256*4+set_id*16+6], codeword_reg8[256*4+set_id*16+6], codeword_reg7[256*4+set_id*16+6], codeword_reg6[256*4+set_id*16+6], codeword_reg5[256*4+set_id*16+6], codeword_reg4[256*4+set_id*16+6], codeword_reg3[256*4+set_id*16+6], codeword_reg2[256*4+set_id*16+6], codeword_reg1[256*4+set_id*16+6], codeword_reg16[256*3+set_id*16+6], codeword_reg15[256*3+set_id*16+6], codeword_reg14[256*3+set_id*16+6], codeword_reg13[256*3+set_id*16+6], codeword_reg12[256*3+set_id*16+6], codeword_reg11[256*3+set_id*16+6], codeword_reg10[256*3+set_id*16+6], codeword_reg9[256*3+set_id*16+6], codeword_reg8[256*3+set_id*16+6], codeword_reg7[256*3+set_id*16+6], codeword_reg6[256*3+set_id*16+6], codeword_reg5[256*3+set_id*16+6], codeword_reg4[256*3+set_id*16+6], codeword_reg3[256*3+set_id*16+6], codeword_reg2[256*3+set_id*16+6], codeword_reg1[256*3+set_id*16+6], codeword_reg16[256*2+set_id*16+6], codeword_reg15[256*2+set_id*16+6], codeword_reg14[256*2+set_id*16+6], codeword_reg13[256*2+set_id*16+6], codeword_reg12[256*2+set_id*16+6], codeword_reg11[256*2+set_id*16+6], codeword_reg10[256*2+set_id*16+6], codeword_reg9[256*2+set_id*16+6], codeword_reg8[256*2+set_id*16+6], codeword_reg7[256*2+set_id*16+6], codeword_reg6[256*2+set_id*16+6], codeword_reg5[256*2+set_id*16+6], codeword_reg4[256*2+set_id*16+6], codeword_reg3[256*2+set_id*16+6], codeword_reg2[256*2+set_id*16+6], codeword_reg1[256*2+set_id*16+6], codeword_reg16[256*1+set_id*16+6], codeword_reg15[256*1+set_id*16+6], codeword_reg14[256*1+set_id*16+6], codeword_reg13[256*1+set_id*16+6], codeword_reg12[256*1+set_id*16+6], codeword_reg11[256*1+set_id*16+6], codeword_reg10[256*1+set_id*16+6], codeword_reg9[256*1+set_id*16+6], codeword_reg8[256*1+set_id*16+6], codeword_reg7[256*1+set_id*16+6], codeword_reg6[256*1+set_id*16+6], codeword_reg5[256*1+set_id*16+6], codeword_reg4[256*1+set_id*16+6], codeword_reg3[256*1+set_id*16+6], codeword_reg2[256*1+set_id*16+6], codeword_reg1[256*1+set_id*16+6], codeword_reg16[256*0+set_id*16+6], codeword_reg15[256*0+set_id*16+6], codeword_reg14[256*0+set_id*16+6], codeword_reg13[256*0+set_id*16+6], codeword_reg12[256*0+set_id*16+6], codeword_reg11[256*0+set_id*16+6], codeword_reg10[256*0+set_id*16+6], codeword_reg9[256*0+set_id*16+6], codeword_reg8[256*0+set_id*16+6], codeword_reg7[256*0+set_id*16+6], codeword_reg6[256*0+set_id*16+6], codeword_reg5[256*0+set_id*16+6], codeword_reg4[256*0+set_id*16+6], codeword_reg3[256*0+set_id*16+6], codeword_reg2[256*0+set_id*16+6], codeword_reg1[256*0+set_id*16+6]};
                            in_bits8  <= {codeword_reg16[256*14+set_id*16+7], codeword_reg15[256*14+set_id*16+7], codeword_reg14[256*14+set_id*16+7], codeword_reg13[256*14+set_id*16+7], codeword_reg12[256*14+set_id*16+7], codeword_reg11[256*14+set_id*16+7], codeword_reg10[256*14+set_id*16+7], codeword_reg9[256*14+set_id*16+7], codeword_reg8[256*14+set_id*16+7], codeword_reg7[256*14+set_id*16+7], codeword_reg6[256*14+set_id*16+7], codeword_reg5[256*14+set_id*16+7], codeword_reg4[256*14+set_id*16+7], codeword_reg3[256*14+set_id*16+7], codeword_reg2[256*14+set_id*16+7], codeword_reg1[256*14+set_id*16+7], codeword_reg16[256*13+set_id*16+7], codeword_reg15[256*13+set_id*16+7], codeword_reg14[256*13+set_id*16+7], codeword_reg13[256*13+set_id*16+7], codeword_reg12[256*13+set_id*16+7], codeword_reg11[256*13+set_id*16+7], codeword_reg10[256*13+set_id*16+7], codeword_reg9[256*13+set_id*16+7], codeword_reg8[256*13+set_id*16+7], codeword_reg7[256*13+set_id*16+7], codeword_reg6[256*13+set_id*16+7], codeword_reg5[256*13+set_id*16+7], codeword_reg4[256*13+set_id*16+7], codeword_reg3[256*13+set_id*16+7], codeword_reg2[256*13+set_id*16+7], codeword_reg1[256*13+set_id*16+7], codeword_reg16[256*12+set_id*16+7], codeword_reg15[256*12+set_id*16+7], codeword_reg14[256*12+set_id*16+7], codeword_reg13[256*12+set_id*16+7], codeword_reg12[256*12+set_id*16+7], codeword_reg11[256*12+set_id*16+7], codeword_reg10[256*12+set_id*16+7], codeword_reg9[256*12+set_id*16+7], codeword_reg8[256*12+set_id*16+7], codeword_reg7[256*12+set_id*16+7], codeword_reg6[256*12+set_id*16+7], codeword_reg5[256*12+set_id*16+7], codeword_reg4[256*12+set_id*16+7], codeword_reg3[256*12+set_id*16+7], codeword_reg2[256*12+set_id*16+7], codeword_reg1[256*12+set_id*16+7], codeword_reg16[256*11+set_id*16+7], codeword_reg15[256*11+set_id*16+7], codeword_reg14[256*11+set_id*16+7], codeword_reg13[256*11+set_id*16+7], codeword_reg12[256*11+set_id*16+7], codeword_reg11[256*11+set_id*16+7], codeword_reg10[256*11+set_id*16+7], codeword_reg9[256*11+set_id*16+7], codeword_reg8[256*11+set_id*16+7], codeword_reg7[256*11+set_id*16+7], codeword_reg6[256*11+set_id*16+7], codeword_reg5[256*11+set_id*16+7], codeword_reg4[256*11+set_id*16+7], codeword_reg3[256*11+set_id*16+7], codeword_reg2[256*11+set_id*16+7], codeword_reg1[256*11+set_id*16+7], codeword_reg16[256*10+set_id*16+7], codeword_reg15[256*10+set_id*16+7], codeword_reg14[256*10+set_id*16+7], codeword_reg13[256*10+set_id*16+7], codeword_reg12[256*10+set_id*16+7], codeword_reg11[256*10+set_id*16+7], codeword_reg10[256*10+set_id*16+7], codeword_reg9[256*10+set_id*16+7], codeword_reg8[256*10+set_id*16+7], codeword_reg7[256*10+set_id*16+7], codeword_reg6[256*10+set_id*16+7], codeword_reg5[256*10+set_id*16+7], codeword_reg4[256*10+set_id*16+7], codeword_reg3[256*10+set_id*16+7], codeword_reg2[256*10+set_id*16+7], codeword_reg1[256*10+set_id*16+7], codeword_reg16[256*9+set_id*16+7], codeword_reg15[256*9+set_id*16+7], codeword_reg14[256*9+set_id*16+7], codeword_reg13[256*9+set_id*16+7], codeword_reg12[256*9+set_id*16+7], codeword_reg11[256*9+set_id*16+7], codeword_reg10[256*9+set_id*16+7], codeword_reg9[256*9+set_id*16+7], codeword_reg8[256*9+set_id*16+7], codeword_reg7[256*9+set_id*16+7], codeword_reg6[256*9+set_id*16+7], codeword_reg5[256*9+set_id*16+7], codeword_reg4[256*9+set_id*16+7], codeword_reg3[256*9+set_id*16+7], codeword_reg2[256*9+set_id*16+7], codeword_reg1[256*9+set_id*16+7], codeword_reg16[256*8+set_id*16+7], codeword_reg15[256*8+set_id*16+7], codeword_reg14[256*8+set_id*16+7], codeword_reg13[256*8+set_id*16+7], codeword_reg12[256*8+set_id*16+7], codeword_reg11[256*8+set_id*16+7], codeword_reg10[256*8+set_id*16+7], codeword_reg9[256*8+set_id*16+7], codeword_reg8[256*8+set_id*16+7], codeword_reg7[256*8+set_id*16+7], codeword_reg6[256*8+set_id*16+7], codeword_reg5[256*8+set_id*16+7], codeword_reg4[256*8+set_id*16+7], codeword_reg3[256*8+set_id*16+7], codeword_reg2[256*8+set_id*16+7], codeword_reg1[256*8+set_id*16+7], codeword_reg16[256*7+set_id*16+7], codeword_reg15[256*7+set_id*16+7], codeword_reg14[256*7+set_id*16+7], codeword_reg13[256*7+set_id*16+7], codeword_reg12[256*7+set_id*16+7], codeword_reg11[256*7+set_id*16+7], codeword_reg10[256*7+set_id*16+7], codeword_reg9[256*7+set_id*16+7], codeword_reg8[256*7+set_id*16+7], codeword_reg7[256*7+set_id*16+7], codeword_reg6[256*7+set_id*16+7], codeword_reg5[256*7+set_id*16+7], codeword_reg4[256*7+set_id*16+7], codeword_reg3[256*7+set_id*16+7], codeword_reg2[256*7+set_id*16+7], codeword_reg1[256*7+set_id*16+7], codeword_reg16[256*6+set_id*16+7], codeword_reg15[256*6+set_id*16+7], codeword_reg14[256*6+set_id*16+7], codeword_reg13[256*6+set_id*16+7], codeword_reg12[256*6+set_id*16+7], codeword_reg11[256*6+set_id*16+7], codeword_reg10[256*6+set_id*16+7], codeword_reg9[256*6+set_id*16+7], codeword_reg8[256*6+set_id*16+7], codeword_reg7[256*6+set_id*16+7], codeword_reg6[256*6+set_id*16+7], codeword_reg5[256*6+set_id*16+7], codeword_reg4[256*6+set_id*16+7], codeword_reg3[256*6+set_id*16+7], codeword_reg2[256*6+set_id*16+7], codeword_reg1[256*6+set_id*16+7], codeword_reg16[256*5+set_id*16+7], codeword_reg15[256*5+set_id*16+7], codeword_reg14[256*5+set_id*16+7], codeword_reg13[256*5+set_id*16+7], codeword_reg12[256*5+set_id*16+7], codeword_reg11[256*5+set_id*16+7], codeword_reg10[256*5+set_id*16+7], codeword_reg9[256*5+set_id*16+7], codeword_reg8[256*5+set_id*16+7], codeword_reg7[256*5+set_id*16+7], codeword_reg6[256*5+set_id*16+7], codeword_reg5[256*5+set_id*16+7], codeword_reg4[256*5+set_id*16+7], codeword_reg3[256*5+set_id*16+7], codeword_reg2[256*5+set_id*16+7], codeword_reg1[256*5+set_id*16+7], codeword_reg16[256*4+set_id*16+7], codeword_reg15[256*4+set_id*16+7], codeword_reg14[256*4+set_id*16+7], codeword_reg13[256*4+set_id*16+7], codeword_reg12[256*4+set_id*16+7], codeword_reg11[256*4+set_id*16+7], codeword_reg10[256*4+set_id*16+7], codeword_reg9[256*4+set_id*16+7], codeword_reg8[256*4+set_id*16+7], codeword_reg7[256*4+set_id*16+7], codeword_reg6[256*4+set_id*16+7], codeword_reg5[256*4+set_id*16+7], codeword_reg4[256*4+set_id*16+7], codeword_reg3[256*4+set_id*16+7], codeword_reg2[256*4+set_id*16+7], codeword_reg1[256*4+set_id*16+7], codeword_reg16[256*3+set_id*16+7], codeword_reg15[256*3+set_id*16+7], codeword_reg14[256*3+set_id*16+7], codeword_reg13[256*3+set_id*16+7], codeword_reg12[256*3+set_id*16+7], codeword_reg11[256*3+set_id*16+7], codeword_reg10[256*3+set_id*16+7], codeword_reg9[256*3+set_id*16+7], codeword_reg8[256*3+set_id*16+7], codeword_reg7[256*3+set_id*16+7], codeword_reg6[256*3+set_id*16+7], codeword_reg5[256*3+set_id*16+7], codeword_reg4[256*3+set_id*16+7], codeword_reg3[256*3+set_id*16+7], codeword_reg2[256*3+set_id*16+7], codeword_reg1[256*3+set_id*16+7], codeword_reg16[256*2+set_id*16+7], codeword_reg15[256*2+set_id*16+7], codeword_reg14[256*2+set_id*16+7], codeword_reg13[256*2+set_id*16+7], codeword_reg12[256*2+set_id*16+7], codeword_reg11[256*2+set_id*16+7], codeword_reg10[256*2+set_id*16+7], codeword_reg9[256*2+set_id*16+7], codeword_reg8[256*2+set_id*16+7], codeword_reg7[256*2+set_id*16+7], codeword_reg6[256*2+set_id*16+7], codeword_reg5[256*2+set_id*16+7], codeword_reg4[256*2+set_id*16+7], codeword_reg3[256*2+set_id*16+7], codeword_reg2[256*2+set_id*16+7], codeword_reg1[256*2+set_id*16+7], codeword_reg16[256*1+set_id*16+7], codeword_reg15[256*1+set_id*16+7], codeword_reg14[256*1+set_id*16+7], codeword_reg13[256*1+set_id*16+7], codeword_reg12[256*1+set_id*16+7], codeword_reg11[256*1+set_id*16+7], codeword_reg10[256*1+set_id*16+7], codeword_reg9[256*1+set_id*16+7], codeword_reg8[256*1+set_id*16+7], codeword_reg7[256*1+set_id*16+7], codeword_reg6[256*1+set_id*16+7], codeword_reg5[256*1+set_id*16+7], codeword_reg4[256*1+set_id*16+7], codeword_reg3[256*1+set_id*16+7], codeword_reg2[256*1+set_id*16+7], codeword_reg1[256*1+set_id*16+7], codeword_reg16[256*0+set_id*16+7], codeword_reg15[256*0+set_id*16+7], codeword_reg14[256*0+set_id*16+7], codeword_reg13[256*0+set_id*16+7], codeword_reg12[256*0+set_id*16+7], codeword_reg11[256*0+set_id*16+7], codeword_reg10[256*0+set_id*16+7], codeword_reg9[256*0+set_id*16+7], codeword_reg8[256*0+set_id*16+7], codeword_reg7[256*0+set_id*16+7], codeword_reg6[256*0+set_id*16+7], codeword_reg5[256*0+set_id*16+7], codeword_reg4[256*0+set_id*16+7], codeword_reg3[256*0+set_id*16+7], codeword_reg2[256*0+set_id*16+7], codeword_reg1[256*0+set_id*16+7]};
                            in_bits9  <= {codeword_reg16[256*14+set_id*16+8], codeword_reg15[256*14+set_id*16+8], codeword_reg14[256*14+set_id*16+8], codeword_reg13[256*14+set_id*16+8], codeword_reg12[256*14+set_id*16+8], codeword_reg11[256*14+set_id*16+8], codeword_reg10[256*14+set_id*16+8], codeword_reg9[256*14+set_id*16+8], codeword_reg8[256*14+set_id*16+8], codeword_reg7[256*14+set_id*16+8], codeword_reg6[256*14+set_id*16+8], codeword_reg5[256*14+set_id*16+8], codeword_reg4[256*14+set_id*16+8], codeword_reg3[256*14+set_id*16+8], codeword_reg2[256*14+set_id*16+8], codeword_reg1[256*14+set_id*16+8], codeword_reg16[256*13+set_id*16+8], codeword_reg15[256*13+set_id*16+8], codeword_reg14[256*13+set_id*16+8], codeword_reg13[256*13+set_id*16+8], codeword_reg12[256*13+set_id*16+8], codeword_reg11[256*13+set_id*16+8], codeword_reg10[256*13+set_id*16+8], codeword_reg9[256*13+set_id*16+8], codeword_reg8[256*13+set_id*16+8], codeword_reg7[256*13+set_id*16+8], codeword_reg6[256*13+set_id*16+8], codeword_reg5[256*13+set_id*16+8], codeword_reg4[256*13+set_id*16+8], codeword_reg3[256*13+set_id*16+8], codeword_reg2[256*13+set_id*16+8], codeword_reg1[256*13+set_id*16+8], codeword_reg16[256*12+set_id*16+8], codeword_reg15[256*12+set_id*16+8], codeword_reg14[256*12+set_id*16+8], codeword_reg13[256*12+set_id*16+8], codeword_reg12[256*12+set_id*16+8], codeword_reg11[256*12+set_id*16+8], codeword_reg10[256*12+set_id*16+8], codeword_reg9[256*12+set_id*16+8], codeword_reg8[256*12+set_id*16+8], codeword_reg7[256*12+set_id*16+8], codeword_reg6[256*12+set_id*16+8], codeword_reg5[256*12+set_id*16+8], codeword_reg4[256*12+set_id*16+8], codeword_reg3[256*12+set_id*16+8], codeword_reg2[256*12+set_id*16+8], codeword_reg1[256*12+set_id*16+8], codeword_reg16[256*11+set_id*16+8], codeword_reg15[256*11+set_id*16+8], codeword_reg14[256*11+set_id*16+8], codeword_reg13[256*11+set_id*16+8], codeword_reg12[256*11+set_id*16+8], codeword_reg11[256*11+set_id*16+8], codeword_reg10[256*11+set_id*16+8], codeword_reg9[256*11+set_id*16+8], codeword_reg8[256*11+set_id*16+8], codeword_reg7[256*11+set_id*16+8], codeword_reg6[256*11+set_id*16+8], codeword_reg5[256*11+set_id*16+8], codeword_reg4[256*11+set_id*16+8], codeword_reg3[256*11+set_id*16+8], codeword_reg2[256*11+set_id*16+8], codeword_reg1[256*11+set_id*16+8], codeword_reg16[256*10+set_id*16+8], codeword_reg15[256*10+set_id*16+8], codeword_reg14[256*10+set_id*16+8], codeword_reg13[256*10+set_id*16+8], codeword_reg12[256*10+set_id*16+8], codeword_reg11[256*10+set_id*16+8], codeword_reg10[256*10+set_id*16+8], codeword_reg9[256*10+set_id*16+8], codeword_reg8[256*10+set_id*16+8], codeword_reg7[256*10+set_id*16+8], codeword_reg6[256*10+set_id*16+8], codeword_reg5[256*10+set_id*16+8], codeword_reg4[256*10+set_id*16+8], codeword_reg3[256*10+set_id*16+8], codeword_reg2[256*10+set_id*16+8], codeword_reg1[256*10+set_id*16+8], codeword_reg16[256*9+set_id*16+8], codeword_reg15[256*9+set_id*16+8], codeword_reg14[256*9+set_id*16+8], codeword_reg13[256*9+set_id*16+8], codeword_reg12[256*9+set_id*16+8], codeword_reg11[256*9+set_id*16+8], codeword_reg10[256*9+set_id*16+8], codeword_reg9[256*9+set_id*16+8], codeword_reg8[256*9+set_id*16+8], codeword_reg7[256*9+set_id*16+8], codeword_reg6[256*9+set_id*16+8], codeword_reg5[256*9+set_id*16+8], codeword_reg4[256*9+set_id*16+8], codeword_reg3[256*9+set_id*16+8], codeword_reg2[256*9+set_id*16+8], codeword_reg1[256*9+set_id*16+8], codeword_reg16[256*8+set_id*16+8], codeword_reg15[256*8+set_id*16+8], codeword_reg14[256*8+set_id*16+8], codeword_reg13[256*8+set_id*16+8], codeword_reg12[256*8+set_id*16+8], codeword_reg11[256*8+set_id*16+8], codeword_reg10[256*8+set_id*16+8], codeword_reg9[256*8+set_id*16+8], codeword_reg8[256*8+set_id*16+8], codeword_reg7[256*8+set_id*16+8], codeword_reg6[256*8+set_id*16+8], codeword_reg5[256*8+set_id*16+8], codeword_reg4[256*8+set_id*16+8], codeword_reg3[256*8+set_id*16+8], codeword_reg2[256*8+set_id*16+8], codeword_reg1[256*8+set_id*16+8], codeword_reg16[256*7+set_id*16+8], codeword_reg15[256*7+set_id*16+8], codeword_reg14[256*7+set_id*16+8], codeword_reg13[256*7+set_id*16+8], codeword_reg12[256*7+set_id*16+8], codeword_reg11[256*7+set_id*16+8], codeword_reg10[256*7+set_id*16+8], codeword_reg9[256*7+set_id*16+8], codeword_reg8[256*7+set_id*16+8], codeword_reg7[256*7+set_id*16+8], codeword_reg6[256*7+set_id*16+8], codeword_reg5[256*7+set_id*16+8], codeword_reg4[256*7+set_id*16+8], codeword_reg3[256*7+set_id*16+8], codeword_reg2[256*7+set_id*16+8], codeword_reg1[256*7+set_id*16+8], codeword_reg16[256*6+set_id*16+8], codeword_reg15[256*6+set_id*16+8], codeword_reg14[256*6+set_id*16+8], codeword_reg13[256*6+set_id*16+8], codeword_reg12[256*6+set_id*16+8], codeword_reg11[256*6+set_id*16+8], codeword_reg10[256*6+set_id*16+8], codeword_reg9[256*6+set_id*16+8], codeword_reg8[256*6+set_id*16+8], codeword_reg7[256*6+set_id*16+8], codeword_reg6[256*6+set_id*16+8], codeword_reg5[256*6+set_id*16+8], codeword_reg4[256*6+set_id*16+8], codeword_reg3[256*6+set_id*16+8], codeword_reg2[256*6+set_id*16+8], codeword_reg1[256*6+set_id*16+8], codeword_reg16[256*5+set_id*16+8], codeword_reg15[256*5+set_id*16+8], codeword_reg14[256*5+set_id*16+8], codeword_reg13[256*5+set_id*16+8], codeword_reg12[256*5+set_id*16+8], codeword_reg11[256*5+set_id*16+8], codeword_reg10[256*5+set_id*16+8], codeword_reg9[256*5+set_id*16+8], codeword_reg8[256*5+set_id*16+8], codeword_reg7[256*5+set_id*16+8], codeword_reg6[256*5+set_id*16+8], codeword_reg5[256*5+set_id*16+8], codeword_reg4[256*5+set_id*16+8], codeword_reg3[256*5+set_id*16+8], codeword_reg2[256*5+set_id*16+8], codeword_reg1[256*5+set_id*16+8], codeword_reg16[256*4+set_id*16+8], codeword_reg15[256*4+set_id*16+8], codeword_reg14[256*4+set_id*16+8], codeword_reg13[256*4+set_id*16+8], codeword_reg12[256*4+set_id*16+8], codeword_reg11[256*4+set_id*16+8], codeword_reg10[256*4+set_id*16+8], codeword_reg9[256*4+set_id*16+8], codeword_reg8[256*4+set_id*16+8], codeword_reg7[256*4+set_id*16+8], codeword_reg6[256*4+set_id*16+8], codeword_reg5[256*4+set_id*16+8], codeword_reg4[256*4+set_id*16+8], codeword_reg3[256*4+set_id*16+8], codeword_reg2[256*4+set_id*16+8], codeword_reg1[256*4+set_id*16+8], codeword_reg16[256*3+set_id*16+8], codeword_reg15[256*3+set_id*16+8], codeword_reg14[256*3+set_id*16+8], codeword_reg13[256*3+set_id*16+8], codeword_reg12[256*3+set_id*16+8], codeword_reg11[256*3+set_id*16+8], codeword_reg10[256*3+set_id*16+8], codeword_reg9[256*3+set_id*16+8], codeword_reg8[256*3+set_id*16+8], codeword_reg7[256*3+set_id*16+8], codeword_reg6[256*3+set_id*16+8], codeword_reg5[256*3+set_id*16+8], codeword_reg4[256*3+set_id*16+8], codeword_reg3[256*3+set_id*16+8], codeword_reg2[256*3+set_id*16+8], codeword_reg1[256*3+set_id*16+8], codeword_reg16[256*2+set_id*16+8], codeword_reg15[256*2+set_id*16+8], codeword_reg14[256*2+set_id*16+8], codeword_reg13[256*2+set_id*16+8], codeword_reg12[256*2+set_id*16+8], codeword_reg11[256*2+set_id*16+8], codeword_reg10[256*2+set_id*16+8], codeword_reg9[256*2+set_id*16+8], codeword_reg8[256*2+set_id*16+8], codeword_reg7[256*2+set_id*16+8], codeword_reg6[256*2+set_id*16+8], codeword_reg5[256*2+set_id*16+8], codeword_reg4[256*2+set_id*16+8], codeword_reg3[256*2+set_id*16+8], codeword_reg2[256*2+set_id*16+8], codeword_reg1[256*2+set_id*16+8], codeword_reg16[256*1+set_id*16+8], codeword_reg15[256*1+set_id*16+8], codeword_reg14[256*1+set_id*16+8], codeword_reg13[256*1+set_id*16+8], codeword_reg12[256*1+set_id*16+8], codeword_reg11[256*1+set_id*16+8], codeword_reg10[256*1+set_id*16+8], codeword_reg9[256*1+set_id*16+8], codeword_reg8[256*1+set_id*16+8], codeword_reg7[256*1+set_id*16+8], codeword_reg6[256*1+set_id*16+8], codeword_reg5[256*1+set_id*16+8], codeword_reg4[256*1+set_id*16+8], codeword_reg3[256*1+set_id*16+8], codeword_reg2[256*1+set_id*16+8], codeword_reg1[256*1+set_id*16+8], codeword_reg16[256*0+set_id*16+8], codeword_reg15[256*0+set_id*16+8], codeword_reg14[256*0+set_id*16+8], codeword_reg13[256*0+set_id*16+8], codeword_reg12[256*0+set_id*16+8], codeword_reg11[256*0+set_id*16+8], codeword_reg10[256*0+set_id*16+8], codeword_reg9[256*0+set_id*16+8], codeword_reg8[256*0+set_id*16+8], codeword_reg7[256*0+set_id*16+8], codeword_reg6[256*0+set_id*16+8], codeword_reg5[256*0+set_id*16+8], codeword_reg4[256*0+set_id*16+8], codeword_reg3[256*0+set_id*16+8], codeword_reg2[256*0+set_id*16+8], codeword_reg1[256*0+set_id*16+8]};
                            in_bits10 <= {codeword_reg16[256*14+set_id*16+9], codeword_reg15[256*14+set_id*16+9], codeword_reg14[256*14+set_id*16+9], codeword_reg13[256*14+set_id*16+9], codeword_reg12[256*14+set_id*16+9], codeword_reg11[256*14+set_id*16+9], codeword_reg10[256*14+set_id*16+9], codeword_reg9[256*14+set_id*16+9], codeword_reg8[256*14+set_id*16+9], codeword_reg7[256*14+set_id*16+9], codeword_reg6[256*14+set_id*16+9], codeword_reg5[256*14+set_id*16+9], codeword_reg4[256*14+set_id*16+9], codeword_reg3[256*14+set_id*16+9], codeword_reg2[256*14+set_id*16+9], codeword_reg1[256*14+set_id*16+9], codeword_reg16[256*13+set_id*16+9], codeword_reg15[256*13+set_id*16+9], codeword_reg14[256*13+set_id*16+9], codeword_reg13[256*13+set_id*16+9], codeword_reg12[256*13+set_id*16+9], codeword_reg11[256*13+set_id*16+9], codeword_reg10[256*13+set_id*16+9], codeword_reg9[256*13+set_id*16+9], codeword_reg8[256*13+set_id*16+9], codeword_reg7[256*13+set_id*16+9], codeword_reg6[256*13+set_id*16+9], codeword_reg5[256*13+set_id*16+9], codeword_reg4[256*13+set_id*16+9], codeword_reg3[256*13+set_id*16+9], codeword_reg2[256*13+set_id*16+9], codeword_reg1[256*13+set_id*16+9], codeword_reg16[256*12+set_id*16+9], codeword_reg15[256*12+set_id*16+9], codeword_reg14[256*12+set_id*16+9], codeword_reg13[256*12+set_id*16+9], codeword_reg12[256*12+set_id*16+9], codeword_reg11[256*12+set_id*16+9], codeword_reg10[256*12+set_id*16+9], codeword_reg9[256*12+set_id*16+9], codeword_reg8[256*12+set_id*16+9], codeword_reg7[256*12+set_id*16+9], codeword_reg6[256*12+set_id*16+9], codeword_reg5[256*12+set_id*16+9], codeword_reg4[256*12+set_id*16+9], codeword_reg3[256*12+set_id*16+9], codeword_reg2[256*12+set_id*16+9], codeword_reg1[256*12+set_id*16+9], codeword_reg16[256*11+set_id*16+9], codeword_reg15[256*11+set_id*16+9], codeword_reg14[256*11+set_id*16+9], codeword_reg13[256*11+set_id*16+9], codeword_reg12[256*11+set_id*16+9], codeword_reg11[256*11+set_id*16+9], codeword_reg10[256*11+set_id*16+9], codeword_reg9[256*11+set_id*16+9], codeword_reg8[256*11+set_id*16+9], codeword_reg7[256*11+set_id*16+9], codeword_reg6[256*11+set_id*16+9], codeword_reg5[256*11+set_id*16+9], codeword_reg4[256*11+set_id*16+9], codeword_reg3[256*11+set_id*16+9], codeword_reg2[256*11+set_id*16+9], codeword_reg1[256*11+set_id*16+9], codeword_reg16[256*10+set_id*16+9], codeword_reg15[256*10+set_id*16+9], codeword_reg14[256*10+set_id*16+9], codeword_reg13[256*10+set_id*16+9], codeword_reg12[256*10+set_id*16+9], codeword_reg11[256*10+set_id*16+9], codeword_reg10[256*10+set_id*16+9], codeword_reg9[256*10+set_id*16+9], codeword_reg8[256*10+set_id*16+9], codeword_reg7[256*10+set_id*16+9], codeword_reg6[256*10+set_id*16+9], codeword_reg5[256*10+set_id*16+9], codeword_reg4[256*10+set_id*16+9], codeword_reg3[256*10+set_id*16+9], codeword_reg2[256*10+set_id*16+9], codeword_reg1[256*10+set_id*16+9], codeword_reg16[256*9+set_id*16+9], codeword_reg15[256*9+set_id*16+9], codeword_reg14[256*9+set_id*16+9], codeword_reg13[256*9+set_id*16+9], codeword_reg12[256*9+set_id*16+9], codeword_reg11[256*9+set_id*16+9], codeword_reg10[256*9+set_id*16+9], codeword_reg9[256*9+set_id*16+9], codeword_reg8[256*9+set_id*16+9], codeword_reg7[256*9+set_id*16+9], codeword_reg6[256*9+set_id*16+9], codeword_reg5[256*9+set_id*16+9], codeword_reg4[256*9+set_id*16+9], codeword_reg3[256*9+set_id*16+9], codeword_reg2[256*9+set_id*16+9], codeword_reg1[256*9+set_id*16+9], codeword_reg16[256*8+set_id*16+9], codeword_reg15[256*8+set_id*16+9], codeword_reg14[256*8+set_id*16+9], codeword_reg13[256*8+set_id*16+9], codeword_reg12[256*8+set_id*16+9], codeword_reg11[256*8+set_id*16+9], codeword_reg10[256*8+set_id*16+9], codeword_reg9[256*8+set_id*16+9], codeword_reg8[256*8+set_id*16+9], codeword_reg7[256*8+set_id*16+9], codeword_reg6[256*8+set_id*16+9], codeword_reg5[256*8+set_id*16+9], codeword_reg4[256*8+set_id*16+9], codeword_reg3[256*8+set_id*16+9], codeword_reg2[256*8+set_id*16+9], codeword_reg1[256*8+set_id*16+9], codeword_reg16[256*7+set_id*16+9], codeword_reg15[256*7+set_id*16+9], codeword_reg14[256*7+set_id*16+9], codeword_reg13[256*7+set_id*16+9], codeword_reg12[256*7+set_id*16+9], codeword_reg11[256*7+set_id*16+9], codeword_reg10[256*7+set_id*16+9], codeword_reg9[256*7+set_id*16+9], codeword_reg8[256*7+set_id*16+9], codeword_reg7[256*7+set_id*16+9], codeword_reg6[256*7+set_id*16+9], codeword_reg5[256*7+set_id*16+9], codeword_reg4[256*7+set_id*16+9], codeword_reg3[256*7+set_id*16+9], codeword_reg2[256*7+set_id*16+9], codeword_reg1[256*7+set_id*16+9], codeword_reg16[256*6+set_id*16+9], codeword_reg15[256*6+set_id*16+9], codeword_reg14[256*6+set_id*16+9], codeword_reg13[256*6+set_id*16+9], codeword_reg12[256*6+set_id*16+9], codeword_reg11[256*6+set_id*16+9], codeword_reg10[256*6+set_id*16+9], codeword_reg9[256*6+set_id*16+9], codeword_reg8[256*6+set_id*16+9], codeword_reg7[256*6+set_id*16+9], codeword_reg6[256*6+set_id*16+9], codeword_reg5[256*6+set_id*16+9], codeword_reg4[256*6+set_id*16+9], codeword_reg3[256*6+set_id*16+9], codeword_reg2[256*6+set_id*16+9], codeword_reg1[256*6+set_id*16+9], codeword_reg16[256*5+set_id*16+9], codeword_reg15[256*5+set_id*16+9], codeword_reg14[256*5+set_id*16+9], codeword_reg13[256*5+set_id*16+9], codeword_reg12[256*5+set_id*16+9], codeword_reg11[256*5+set_id*16+9], codeword_reg10[256*5+set_id*16+9], codeword_reg9[256*5+set_id*16+9], codeword_reg8[256*5+set_id*16+9], codeword_reg7[256*5+set_id*16+9], codeword_reg6[256*5+set_id*16+9], codeword_reg5[256*5+set_id*16+9], codeword_reg4[256*5+set_id*16+9], codeword_reg3[256*5+set_id*16+9], codeword_reg2[256*5+set_id*16+9], codeword_reg1[256*5+set_id*16+9], codeword_reg16[256*4+set_id*16+9], codeword_reg15[256*4+set_id*16+9], codeword_reg14[256*4+set_id*16+9], codeword_reg13[256*4+set_id*16+9], codeword_reg12[256*4+set_id*16+9], codeword_reg11[256*4+set_id*16+9], codeword_reg10[256*4+set_id*16+9], codeword_reg9[256*4+set_id*16+9], codeword_reg8[256*4+set_id*16+9], codeword_reg7[256*4+set_id*16+9], codeword_reg6[256*4+set_id*16+9], codeword_reg5[256*4+set_id*16+9], codeword_reg4[256*4+set_id*16+9], codeword_reg3[256*4+set_id*16+9], codeword_reg2[256*4+set_id*16+9], codeword_reg1[256*4+set_id*16+9], codeword_reg16[256*3+set_id*16+9], codeword_reg15[256*3+set_id*16+9], codeword_reg14[256*3+set_id*16+9], codeword_reg13[256*3+set_id*16+9], codeword_reg12[256*3+set_id*16+9], codeword_reg11[256*3+set_id*16+9], codeword_reg10[256*3+set_id*16+9], codeword_reg9[256*3+set_id*16+9], codeword_reg8[256*3+set_id*16+9], codeword_reg7[256*3+set_id*16+9], codeword_reg6[256*3+set_id*16+9], codeword_reg5[256*3+set_id*16+9], codeword_reg4[256*3+set_id*16+9], codeword_reg3[256*3+set_id*16+9], codeword_reg2[256*3+set_id*16+9], codeword_reg1[256*3+set_id*16+9], codeword_reg16[256*2+set_id*16+9], codeword_reg15[256*2+set_id*16+9], codeword_reg14[256*2+set_id*16+9], codeword_reg13[256*2+set_id*16+9], codeword_reg12[256*2+set_id*16+9], codeword_reg11[256*2+set_id*16+9], codeword_reg10[256*2+set_id*16+9], codeword_reg9[256*2+set_id*16+9], codeword_reg8[256*2+set_id*16+9], codeword_reg7[256*2+set_id*16+9], codeword_reg6[256*2+set_id*16+9], codeword_reg5[256*2+set_id*16+9], codeword_reg4[256*2+set_id*16+9], codeword_reg3[256*2+set_id*16+9], codeword_reg2[256*2+set_id*16+9], codeword_reg1[256*2+set_id*16+9], codeword_reg16[256*1+set_id*16+9], codeword_reg15[256*1+set_id*16+9], codeword_reg14[256*1+set_id*16+9], codeword_reg13[256*1+set_id*16+9], codeword_reg12[256*1+set_id*16+9], codeword_reg11[256*1+set_id*16+9], codeword_reg10[256*1+set_id*16+9], codeword_reg9[256*1+set_id*16+9], codeword_reg8[256*1+set_id*16+9], codeword_reg7[256*1+set_id*16+9], codeword_reg6[256*1+set_id*16+9], codeword_reg5[256*1+set_id*16+9], codeword_reg4[256*1+set_id*16+9], codeword_reg3[256*1+set_id*16+9], codeword_reg2[256*1+set_id*16+9], codeword_reg1[256*1+set_id*16+9], codeword_reg16[256*0+set_id*16+9], codeword_reg15[256*0+set_id*16+9], codeword_reg14[256*0+set_id*16+9], codeword_reg13[256*0+set_id*16+9], codeword_reg12[256*0+set_id*16+9], codeword_reg11[256*0+set_id*16+9], codeword_reg10[256*0+set_id*16+9], codeword_reg9[256*0+set_id*16+9], codeword_reg8[256*0+set_id*16+9], codeword_reg7[256*0+set_id*16+9], codeword_reg6[256*0+set_id*16+9], codeword_reg5[256*0+set_id*16+9], codeword_reg4[256*0+set_id*16+9], codeword_reg3[256*0+set_id*16+9], codeword_reg2[256*0+set_id*16+9], codeword_reg1[256*0+set_id*16+9]};
                            in_bits11 <= {codeword_reg16[256*14+set_id*16+10], codeword_reg15[256*14+set_id*16+10], codeword_reg14[256*14+set_id*16+10], codeword_reg13[256*14+set_id*16+10], codeword_reg12[256*14+set_id*16+10], codeword_reg11[256*14+set_id*16+10], codeword_reg10[256*14+set_id*16+10], codeword_reg9[256*14+set_id*16+10], codeword_reg8[256*14+set_id*16+10], codeword_reg7[256*14+set_id*16+10], codeword_reg6[256*14+set_id*16+10], codeword_reg5[256*14+set_id*16+10], codeword_reg4[256*14+set_id*16+10], codeword_reg3[256*14+set_id*16+10], codeword_reg2[256*14+set_id*16+10], codeword_reg1[256*14+set_id*16+10], codeword_reg16[256*13+set_id*16+10], codeword_reg15[256*13+set_id*16+10], codeword_reg14[256*13+set_id*16+10], codeword_reg13[256*13+set_id*16+10], codeword_reg12[256*13+set_id*16+10], codeword_reg11[256*13+set_id*16+10], codeword_reg10[256*13+set_id*16+10], codeword_reg9[256*13+set_id*16+10], codeword_reg8[256*13+set_id*16+10], codeword_reg7[256*13+set_id*16+10], codeword_reg6[256*13+set_id*16+10], codeword_reg5[256*13+set_id*16+10], codeword_reg4[256*13+set_id*16+10], codeword_reg3[256*13+set_id*16+10], codeword_reg2[256*13+set_id*16+10], codeword_reg1[256*13+set_id*16+10], codeword_reg16[256*12+set_id*16+10], codeword_reg15[256*12+set_id*16+10], codeword_reg14[256*12+set_id*16+10], codeword_reg13[256*12+set_id*16+10], codeword_reg12[256*12+set_id*16+10], codeword_reg11[256*12+set_id*16+10], codeword_reg10[256*12+set_id*16+10], codeword_reg9[256*12+set_id*16+10], codeword_reg8[256*12+set_id*16+10], codeword_reg7[256*12+set_id*16+10], codeword_reg6[256*12+set_id*16+10], codeword_reg5[256*12+set_id*16+10], codeword_reg4[256*12+set_id*16+10], codeword_reg3[256*12+set_id*16+10], codeword_reg2[256*12+set_id*16+10], codeword_reg1[256*12+set_id*16+10], codeword_reg16[256*11+set_id*16+10], codeword_reg15[256*11+set_id*16+10], codeword_reg14[256*11+set_id*16+10], codeword_reg13[256*11+set_id*16+10], codeword_reg12[256*11+set_id*16+10], codeword_reg11[256*11+set_id*16+10], codeword_reg10[256*11+set_id*16+10], codeword_reg9[256*11+set_id*16+10], codeword_reg8[256*11+set_id*16+10], codeword_reg7[256*11+set_id*16+10], codeword_reg6[256*11+set_id*16+10], codeword_reg5[256*11+set_id*16+10], codeword_reg4[256*11+set_id*16+10], codeword_reg3[256*11+set_id*16+10], codeword_reg2[256*11+set_id*16+10], codeword_reg1[256*11+set_id*16+10], codeword_reg16[256*10+set_id*16+10], codeword_reg15[256*10+set_id*16+10], codeword_reg14[256*10+set_id*16+10], codeword_reg13[256*10+set_id*16+10], codeword_reg12[256*10+set_id*16+10], codeword_reg11[256*10+set_id*16+10], codeword_reg10[256*10+set_id*16+10], codeword_reg9[256*10+set_id*16+10], codeword_reg8[256*10+set_id*16+10], codeword_reg7[256*10+set_id*16+10], codeword_reg6[256*10+set_id*16+10], codeword_reg5[256*10+set_id*16+10], codeword_reg4[256*10+set_id*16+10], codeword_reg3[256*10+set_id*16+10], codeword_reg2[256*10+set_id*16+10], codeword_reg1[256*10+set_id*16+10], codeword_reg16[256*9+set_id*16+10], codeword_reg15[256*9+set_id*16+10], codeword_reg14[256*9+set_id*16+10], codeword_reg13[256*9+set_id*16+10], codeword_reg12[256*9+set_id*16+10], codeword_reg11[256*9+set_id*16+10], codeword_reg10[256*9+set_id*16+10], codeword_reg9[256*9+set_id*16+10], codeword_reg8[256*9+set_id*16+10], codeword_reg7[256*9+set_id*16+10], codeword_reg6[256*9+set_id*16+10], codeword_reg5[256*9+set_id*16+10], codeword_reg4[256*9+set_id*16+10], codeword_reg3[256*9+set_id*16+10], codeword_reg2[256*9+set_id*16+10], codeword_reg1[256*9+set_id*16+10], codeword_reg16[256*8+set_id*16+10], codeword_reg15[256*8+set_id*16+10], codeword_reg14[256*8+set_id*16+10], codeword_reg13[256*8+set_id*16+10], codeword_reg12[256*8+set_id*16+10], codeword_reg11[256*8+set_id*16+10], codeword_reg10[256*8+set_id*16+10], codeword_reg9[256*8+set_id*16+10], codeword_reg8[256*8+set_id*16+10], codeword_reg7[256*8+set_id*16+10], codeword_reg6[256*8+set_id*16+10], codeword_reg5[256*8+set_id*16+10], codeword_reg4[256*8+set_id*16+10], codeword_reg3[256*8+set_id*16+10], codeword_reg2[256*8+set_id*16+10], codeword_reg1[256*8+set_id*16+10], codeword_reg16[256*7+set_id*16+10], codeword_reg15[256*7+set_id*16+10], codeword_reg14[256*7+set_id*16+10], codeword_reg13[256*7+set_id*16+10], codeword_reg12[256*7+set_id*16+10], codeword_reg11[256*7+set_id*16+10], codeword_reg10[256*7+set_id*16+10], codeword_reg9[256*7+set_id*16+10], codeword_reg8[256*7+set_id*16+10], codeword_reg7[256*7+set_id*16+10], codeword_reg6[256*7+set_id*16+10], codeword_reg5[256*7+set_id*16+10], codeword_reg4[256*7+set_id*16+10], codeword_reg3[256*7+set_id*16+10], codeword_reg2[256*7+set_id*16+10], codeword_reg1[256*7+set_id*16+10], codeword_reg16[256*6+set_id*16+10], codeword_reg15[256*6+set_id*16+10], codeword_reg14[256*6+set_id*16+10], codeword_reg13[256*6+set_id*16+10], codeword_reg12[256*6+set_id*16+10], codeword_reg11[256*6+set_id*16+10], codeword_reg10[256*6+set_id*16+10], codeword_reg9[256*6+set_id*16+10], codeword_reg8[256*6+set_id*16+10], codeword_reg7[256*6+set_id*16+10], codeword_reg6[256*6+set_id*16+10], codeword_reg5[256*6+set_id*16+10], codeword_reg4[256*6+set_id*16+10], codeword_reg3[256*6+set_id*16+10], codeword_reg2[256*6+set_id*16+10], codeword_reg1[256*6+set_id*16+10], codeword_reg16[256*5+set_id*16+10], codeword_reg15[256*5+set_id*16+10], codeword_reg14[256*5+set_id*16+10], codeword_reg13[256*5+set_id*16+10], codeword_reg12[256*5+set_id*16+10], codeword_reg11[256*5+set_id*16+10], codeword_reg10[256*5+set_id*16+10], codeword_reg9[256*5+set_id*16+10], codeword_reg8[256*5+set_id*16+10], codeword_reg7[256*5+set_id*16+10], codeword_reg6[256*5+set_id*16+10], codeword_reg5[256*5+set_id*16+10], codeword_reg4[256*5+set_id*16+10], codeword_reg3[256*5+set_id*16+10], codeword_reg2[256*5+set_id*16+10], codeword_reg1[256*5+set_id*16+10], codeword_reg16[256*4+set_id*16+10], codeword_reg15[256*4+set_id*16+10], codeword_reg14[256*4+set_id*16+10], codeword_reg13[256*4+set_id*16+10], codeword_reg12[256*4+set_id*16+10], codeword_reg11[256*4+set_id*16+10], codeword_reg10[256*4+set_id*16+10], codeword_reg9[256*4+set_id*16+10], codeword_reg8[256*4+set_id*16+10], codeword_reg7[256*4+set_id*16+10], codeword_reg6[256*4+set_id*16+10], codeword_reg5[256*4+set_id*16+10], codeword_reg4[256*4+set_id*16+10], codeword_reg3[256*4+set_id*16+10], codeword_reg2[256*4+set_id*16+10], codeword_reg1[256*4+set_id*16+10], codeword_reg16[256*3+set_id*16+10], codeword_reg15[256*3+set_id*16+10], codeword_reg14[256*3+set_id*16+10], codeword_reg13[256*3+set_id*16+10], codeword_reg12[256*3+set_id*16+10], codeword_reg11[256*3+set_id*16+10], codeword_reg10[256*3+set_id*16+10], codeword_reg9[256*3+set_id*16+10], codeword_reg8[256*3+set_id*16+10], codeword_reg7[256*3+set_id*16+10], codeword_reg6[256*3+set_id*16+10], codeword_reg5[256*3+set_id*16+10], codeword_reg4[256*3+set_id*16+10], codeword_reg3[256*3+set_id*16+10], codeword_reg2[256*3+set_id*16+10], codeword_reg1[256*3+set_id*16+10], codeword_reg16[256*2+set_id*16+10], codeword_reg15[256*2+set_id*16+10], codeword_reg14[256*2+set_id*16+10], codeword_reg13[256*2+set_id*16+10], codeword_reg12[256*2+set_id*16+10], codeword_reg11[256*2+set_id*16+10], codeword_reg10[256*2+set_id*16+10], codeword_reg9[256*2+set_id*16+10], codeword_reg8[256*2+set_id*16+10], codeword_reg7[256*2+set_id*16+10], codeword_reg6[256*2+set_id*16+10], codeword_reg5[256*2+set_id*16+10], codeword_reg4[256*2+set_id*16+10], codeword_reg3[256*2+set_id*16+10], codeword_reg2[256*2+set_id*16+10], codeword_reg1[256*2+set_id*16+10], codeword_reg16[256*1+set_id*16+10], codeword_reg15[256*1+set_id*16+10], codeword_reg14[256*1+set_id*16+10], codeword_reg13[256*1+set_id*16+10], codeword_reg12[256*1+set_id*16+10], codeword_reg11[256*1+set_id*16+10], codeword_reg10[256*1+set_id*16+10], codeword_reg9[256*1+set_id*16+10], codeword_reg8[256*1+set_id*16+10], codeword_reg7[256*1+set_id*16+10], codeword_reg6[256*1+set_id*16+10], codeword_reg5[256*1+set_id*16+10], codeword_reg4[256*1+set_id*16+10], codeword_reg3[256*1+set_id*16+10], codeword_reg2[256*1+set_id*16+10], codeword_reg1[256*1+set_id*16+10], codeword_reg16[256*0+set_id*16+10], codeword_reg15[256*0+set_id*16+10], codeword_reg14[256*0+set_id*16+10], codeword_reg13[256*0+set_id*16+10], codeword_reg12[256*0+set_id*16+10], codeword_reg11[256*0+set_id*16+10], codeword_reg10[256*0+set_id*16+10], codeword_reg9[256*0+set_id*16+10], codeword_reg8[256*0+set_id*16+10], codeword_reg7[256*0+set_id*16+10], codeword_reg6[256*0+set_id*16+10], codeword_reg5[256*0+set_id*16+10], codeword_reg4[256*0+set_id*16+10], codeword_reg3[256*0+set_id*16+10], codeword_reg2[256*0+set_id*16+10], codeword_reg1[256*0+set_id*16+10]};
                            in_bits12 <= {codeword_reg16[256*14+set_id*16+11], codeword_reg15[256*14+set_id*16+11], codeword_reg14[256*14+set_id*16+11], codeword_reg13[256*14+set_id*16+11], codeword_reg12[256*14+set_id*16+11], codeword_reg11[256*14+set_id*16+11], codeword_reg10[256*14+set_id*16+11], codeword_reg9[256*14+set_id*16+11], codeword_reg8[256*14+set_id*16+11], codeword_reg7[256*14+set_id*16+11], codeword_reg6[256*14+set_id*16+11], codeword_reg5[256*14+set_id*16+11], codeword_reg4[256*14+set_id*16+11], codeword_reg3[256*14+set_id*16+11], codeword_reg2[256*14+set_id*16+11], codeword_reg1[256*14+set_id*16+11], codeword_reg16[256*13+set_id*16+11], codeword_reg15[256*13+set_id*16+11], codeword_reg14[256*13+set_id*16+11], codeword_reg13[256*13+set_id*16+11], codeword_reg12[256*13+set_id*16+11], codeword_reg11[256*13+set_id*16+11], codeword_reg10[256*13+set_id*16+11], codeword_reg9[256*13+set_id*16+11], codeword_reg8[256*13+set_id*16+11], codeword_reg7[256*13+set_id*16+11], codeword_reg6[256*13+set_id*16+11], codeword_reg5[256*13+set_id*16+11], codeword_reg4[256*13+set_id*16+11], codeword_reg3[256*13+set_id*16+11], codeword_reg2[256*13+set_id*16+11], codeword_reg1[256*13+set_id*16+11], codeword_reg16[256*12+set_id*16+11], codeword_reg15[256*12+set_id*16+11], codeword_reg14[256*12+set_id*16+11], codeword_reg13[256*12+set_id*16+11], codeword_reg12[256*12+set_id*16+11], codeword_reg11[256*12+set_id*16+11], codeword_reg10[256*12+set_id*16+11], codeword_reg9[256*12+set_id*16+11], codeword_reg8[256*12+set_id*16+11], codeword_reg7[256*12+set_id*16+11], codeword_reg6[256*12+set_id*16+11], codeword_reg5[256*12+set_id*16+11], codeword_reg4[256*12+set_id*16+11], codeword_reg3[256*12+set_id*16+11], codeword_reg2[256*12+set_id*16+11], codeword_reg1[256*12+set_id*16+11], codeword_reg16[256*11+set_id*16+11], codeword_reg15[256*11+set_id*16+11], codeword_reg14[256*11+set_id*16+11], codeword_reg13[256*11+set_id*16+11], codeword_reg12[256*11+set_id*16+11], codeword_reg11[256*11+set_id*16+11], codeword_reg10[256*11+set_id*16+11], codeword_reg9[256*11+set_id*16+11], codeword_reg8[256*11+set_id*16+11], codeword_reg7[256*11+set_id*16+11], codeword_reg6[256*11+set_id*16+11], codeword_reg5[256*11+set_id*16+11], codeword_reg4[256*11+set_id*16+11], codeword_reg3[256*11+set_id*16+11], codeword_reg2[256*11+set_id*16+11], codeword_reg1[256*11+set_id*16+11], codeword_reg16[256*10+set_id*16+11], codeword_reg15[256*10+set_id*16+11], codeword_reg14[256*10+set_id*16+11], codeword_reg13[256*10+set_id*16+11], codeword_reg12[256*10+set_id*16+11], codeword_reg11[256*10+set_id*16+11], codeword_reg10[256*10+set_id*16+11], codeword_reg9[256*10+set_id*16+11], codeword_reg8[256*10+set_id*16+11], codeword_reg7[256*10+set_id*16+11], codeword_reg6[256*10+set_id*16+11], codeword_reg5[256*10+set_id*16+11], codeword_reg4[256*10+set_id*16+11], codeword_reg3[256*10+set_id*16+11], codeword_reg2[256*10+set_id*16+11], codeword_reg1[256*10+set_id*16+11], codeword_reg16[256*9+set_id*16+11], codeword_reg15[256*9+set_id*16+11], codeword_reg14[256*9+set_id*16+11], codeword_reg13[256*9+set_id*16+11], codeword_reg12[256*9+set_id*16+11], codeword_reg11[256*9+set_id*16+11], codeword_reg10[256*9+set_id*16+11], codeword_reg9[256*9+set_id*16+11], codeword_reg8[256*9+set_id*16+11], codeword_reg7[256*9+set_id*16+11], codeword_reg6[256*9+set_id*16+11], codeword_reg5[256*9+set_id*16+11], codeword_reg4[256*9+set_id*16+11], codeword_reg3[256*9+set_id*16+11], codeword_reg2[256*9+set_id*16+11], codeword_reg1[256*9+set_id*16+11], codeword_reg16[256*8+set_id*16+11], codeword_reg15[256*8+set_id*16+11], codeword_reg14[256*8+set_id*16+11], codeword_reg13[256*8+set_id*16+11], codeword_reg12[256*8+set_id*16+11], codeword_reg11[256*8+set_id*16+11], codeword_reg10[256*8+set_id*16+11], codeword_reg9[256*8+set_id*16+11], codeword_reg8[256*8+set_id*16+11], codeword_reg7[256*8+set_id*16+11], codeword_reg6[256*8+set_id*16+11], codeword_reg5[256*8+set_id*16+11], codeword_reg4[256*8+set_id*16+11], codeword_reg3[256*8+set_id*16+11], codeword_reg2[256*8+set_id*16+11], codeword_reg1[256*8+set_id*16+11], codeword_reg16[256*7+set_id*16+11], codeword_reg15[256*7+set_id*16+11], codeword_reg14[256*7+set_id*16+11], codeword_reg13[256*7+set_id*16+11], codeword_reg12[256*7+set_id*16+11], codeword_reg11[256*7+set_id*16+11], codeword_reg10[256*7+set_id*16+11], codeword_reg9[256*7+set_id*16+11], codeword_reg8[256*7+set_id*16+11], codeword_reg7[256*7+set_id*16+11], codeword_reg6[256*7+set_id*16+11], codeword_reg5[256*7+set_id*16+11], codeword_reg4[256*7+set_id*16+11], codeword_reg3[256*7+set_id*16+11], codeword_reg2[256*7+set_id*16+11], codeword_reg1[256*7+set_id*16+11], codeword_reg16[256*6+set_id*16+11], codeword_reg15[256*6+set_id*16+11], codeword_reg14[256*6+set_id*16+11], codeword_reg13[256*6+set_id*16+11], codeword_reg12[256*6+set_id*16+11], codeword_reg11[256*6+set_id*16+11], codeword_reg10[256*6+set_id*16+11], codeword_reg9[256*6+set_id*16+11], codeword_reg8[256*6+set_id*16+11], codeword_reg7[256*6+set_id*16+11], codeword_reg6[256*6+set_id*16+11], codeword_reg5[256*6+set_id*16+11], codeword_reg4[256*6+set_id*16+11], codeword_reg3[256*6+set_id*16+11], codeword_reg2[256*6+set_id*16+11], codeword_reg1[256*6+set_id*16+11], codeword_reg16[256*5+set_id*16+11], codeword_reg15[256*5+set_id*16+11], codeword_reg14[256*5+set_id*16+11], codeword_reg13[256*5+set_id*16+11], codeword_reg12[256*5+set_id*16+11], codeword_reg11[256*5+set_id*16+11], codeword_reg10[256*5+set_id*16+11], codeword_reg9[256*5+set_id*16+11], codeword_reg8[256*5+set_id*16+11], codeword_reg7[256*5+set_id*16+11], codeword_reg6[256*5+set_id*16+11], codeword_reg5[256*5+set_id*16+11], codeword_reg4[256*5+set_id*16+11], codeword_reg3[256*5+set_id*16+11], codeword_reg2[256*5+set_id*16+11], codeword_reg1[256*5+set_id*16+11], codeword_reg16[256*4+set_id*16+11], codeword_reg15[256*4+set_id*16+11], codeword_reg14[256*4+set_id*16+11], codeword_reg13[256*4+set_id*16+11], codeword_reg12[256*4+set_id*16+11], codeword_reg11[256*4+set_id*16+11], codeword_reg10[256*4+set_id*16+11], codeword_reg9[256*4+set_id*16+11], codeword_reg8[256*4+set_id*16+11], codeword_reg7[256*4+set_id*16+11], codeword_reg6[256*4+set_id*16+11], codeword_reg5[256*4+set_id*16+11], codeword_reg4[256*4+set_id*16+11], codeword_reg3[256*4+set_id*16+11], codeword_reg2[256*4+set_id*16+11], codeword_reg1[256*4+set_id*16+11], codeword_reg16[256*3+set_id*16+11], codeword_reg15[256*3+set_id*16+11], codeword_reg14[256*3+set_id*16+11], codeword_reg13[256*3+set_id*16+11], codeword_reg12[256*3+set_id*16+11], codeword_reg11[256*3+set_id*16+11], codeword_reg10[256*3+set_id*16+11], codeword_reg9[256*3+set_id*16+11], codeword_reg8[256*3+set_id*16+11], codeword_reg7[256*3+set_id*16+11], codeword_reg6[256*3+set_id*16+11], codeword_reg5[256*3+set_id*16+11], codeword_reg4[256*3+set_id*16+11], codeword_reg3[256*3+set_id*16+11], codeword_reg2[256*3+set_id*16+11], codeword_reg1[256*3+set_id*16+11], codeword_reg16[256*2+set_id*16+11], codeword_reg15[256*2+set_id*16+11], codeword_reg14[256*2+set_id*16+11], codeword_reg13[256*2+set_id*16+11], codeword_reg12[256*2+set_id*16+11], codeword_reg11[256*2+set_id*16+11], codeword_reg10[256*2+set_id*16+11], codeword_reg9[256*2+set_id*16+11], codeword_reg8[256*2+set_id*16+11], codeword_reg7[256*2+set_id*16+11], codeword_reg6[256*2+set_id*16+11], codeword_reg5[256*2+set_id*16+11], codeword_reg4[256*2+set_id*16+11], codeword_reg3[256*2+set_id*16+11], codeword_reg2[256*2+set_id*16+11], codeword_reg1[256*2+set_id*16+11], codeword_reg16[256*1+set_id*16+11], codeword_reg15[256*1+set_id*16+11], codeword_reg14[256*1+set_id*16+11], codeword_reg13[256*1+set_id*16+11], codeword_reg12[256*1+set_id*16+11], codeword_reg11[256*1+set_id*16+11], codeword_reg10[256*1+set_id*16+11], codeword_reg9[256*1+set_id*16+11], codeword_reg8[256*1+set_id*16+11], codeword_reg7[256*1+set_id*16+11], codeword_reg6[256*1+set_id*16+11], codeword_reg5[256*1+set_id*16+11], codeword_reg4[256*1+set_id*16+11], codeword_reg3[256*1+set_id*16+11], codeword_reg2[256*1+set_id*16+11], codeword_reg1[256*1+set_id*16+11], codeword_reg16[256*0+set_id*16+11], codeword_reg15[256*0+set_id*16+11], codeword_reg14[256*0+set_id*16+11], codeword_reg13[256*0+set_id*16+11], codeword_reg12[256*0+set_id*16+11], codeword_reg11[256*0+set_id*16+11], codeword_reg10[256*0+set_id*16+11], codeword_reg9[256*0+set_id*16+11], codeword_reg8[256*0+set_id*16+11], codeword_reg7[256*0+set_id*16+11], codeword_reg6[256*0+set_id*16+11], codeword_reg5[256*0+set_id*16+11], codeword_reg4[256*0+set_id*16+11], codeword_reg3[256*0+set_id*16+11], codeword_reg2[256*0+set_id*16+11], codeword_reg1[256*0+set_id*16+11]};
                            in_bits13 <= {codeword_reg16[256*14+set_id*16+12], codeword_reg15[256*14+set_id*16+12], codeword_reg14[256*14+set_id*16+12], codeword_reg13[256*14+set_id*16+12], codeword_reg12[256*14+set_id*16+12], codeword_reg11[256*14+set_id*16+12], codeword_reg10[256*14+set_id*16+12], codeword_reg9[256*14+set_id*16+12], codeword_reg8[256*14+set_id*16+12], codeword_reg7[256*14+set_id*16+12], codeword_reg6[256*14+set_id*16+12], codeword_reg5[256*14+set_id*16+12], codeword_reg4[256*14+set_id*16+12], codeword_reg3[256*14+set_id*16+12], codeword_reg2[256*14+set_id*16+12], codeword_reg1[256*14+set_id*16+12], codeword_reg16[256*13+set_id*16+12], codeword_reg15[256*13+set_id*16+12], codeword_reg14[256*13+set_id*16+12], codeword_reg13[256*13+set_id*16+12], codeword_reg12[256*13+set_id*16+12], codeword_reg11[256*13+set_id*16+12], codeword_reg10[256*13+set_id*16+12], codeword_reg9[256*13+set_id*16+12], codeword_reg8[256*13+set_id*16+12], codeword_reg7[256*13+set_id*16+12], codeword_reg6[256*13+set_id*16+12], codeword_reg5[256*13+set_id*16+12], codeword_reg4[256*13+set_id*16+12], codeword_reg3[256*13+set_id*16+12], codeword_reg2[256*13+set_id*16+12], codeword_reg1[256*13+set_id*16+12], codeword_reg16[256*12+set_id*16+12], codeword_reg15[256*12+set_id*16+12], codeword_reg14[256*12+set_id*16+12], codeword_reg13[256*12+set_id*16+12], codeword_reg12[256*12+set_id*16+12], codeword_reg11[256*12+set_id*16+12], codeword_reg10[256*12+set_id*16+12], codeword_reg9[256*12+set_id*16+12], codeword_reg8[256*12+set_id*16+12], codeword_reg7[256*12+set_id*16+12], codeword_reg6[256*12+set_id*16+12], codeword_reg5[256*12+set_id*16+12], codeword_reg4[256*12+set_id*16+12], codeword_reg3[256*12+set_id*16+12], codeword_reg2[256*12+set_id*16+12], codeword_reg1[256*12+set_id*16+12], codeword_reg16[256*11+set_id*16+12], codeword_reg15[256*11+set_id*16+12], codeword_reg14[256*11+set_id*16+12], codeword_reg13[256*11+set_id*16+12], codeword_reg12[256*11+set_id*16+12], codeword_reg11[256*11+set_id*16+12], codeword_reg10[256*11+set_id*16+12], codeword_reg9[256*11+set_id*16+12], codeword_reg8[256*11+set_id*16+12], codeword_reg7[256*11+set_id*16+12], codeword_reg6[256*11+set_id*16+12], codeword_reg5[256*11+set_id*16+12], codeword_reg4[256*11+set_id*16+12], codeword_reg3[256*11+set_id*16+12], codeword_reg2[256*11+set_id*16+12], codeword_reg1[256*11+set_id*16+12], codeword_reg16[256*10+set_id*16+12], codeword_reg15[256*10+set_id*16+12], codeword_reg14[256*10+set_id*16+12], codeword_reg13[256*10+set_id*16+12], codeword_reg12[256*10+set_id*16+12], codeword_reg11[256*10+set_id*16+12], codeword_reg10[256*10+set_id*16+12], codeword_reg9[256*10+set_id*16+12], codeword_reg8[256*10+set_id*16+12], codeword_reg7[256*10+set_id*16+12], codeword_reg6[256*10+set_id*16+12], codeword_reg5[256*10+set_id*16+12], codeword_reg4[256*10+set_id*16+12], codeword_reg3[256*10+set_id*16+12], codeword_reg2[256*10+set_id*16+12], codeword_reg1[256*10+set_id*16+12], codeword_reg16[256*9+set_id*16+12], codeword_reg15[256*9+set_id*16+12], codeword_reg14[256*9+set_id*16+12], codeword_reg13[256*9+set_id*16+12], codeword_reg12[256*9+set_id*16+12], codeword_reg11[256*9+set_id*16+12], codeword_reg10[256*9+set_id*16+12], codeword_reg9[256*9+set_id*16+12], codeword_reg8[256*9+set_id*16+12], codeword_reg7[256*9+set_id*16+12], codeword_reg6[256*9+set_id*16+12], codeword_reg5[256*9+set_id*16+12], codeword_reg4[256*9+set_id*16+12], codeword_reg3[256*9+set_id*16+12], codeword_reg2[256*9+set_id*16+12], codeword_reg1[256*9+set_id*16+12], codeword_reg16[256*8+set_id*16+12], codeword_reg15[256*8+set_id*16+12], codeword_reg14[256*8+set_id*16+12], codeword_reg13[256*8+set_id*16+12], codeword_reg12[256*8+set_id*16+12], codeword_reg11[256*8+set_id*16+12], codeword_reg10[256*8+set_id*16+12], codeword_reg9[256*8+set_id*16+12], codeword_reg8[256*8+set_id*16+12], codeword_reg7[256*8+set_id*16+12], codeword_reg6[256*8+set_id*16+12], codeword_reg5[256*8+set_id*16+12], codeword_reg4[256*8+set_id*16+12], codeword_reg3[256*8+set_id*16+12], codeword_reg2[256*8+set_id*16+12], codeword_reg1[256*8+set_id*16+12], codeword_reg16[256*7+set_id*16+12], codeword_reg15[256*7+set_id*16+12], codeword_reg14[256*7+set_id*16+12], codeword_reg13[256*7+set_id*16+12], codeword_reg12[256*7+set_id*16+12], codeword_reg11[256*7+set_id*16+12], codeword_reg10[256*7+set_id*16+12], codeword_reg9[256*7+set_id*16+12], codeword_reg8[256*7+set_id*16+12], codeword_reg7[256*7+set_id*16+12], codeword_reg6[256*7+set_id*16+12], codeword_reg5[256*7+set_id*16+12], codeword_reg4[256*7+set_id*16+12], codeword_reg3[256*7+set_id*16+12], codeword_reg2[256*7+set_id*16+12], codeword_reg1[256*7+set_id*16+12], codeword_reg16[256*6+set_id*16+12], codeword_reg15[256*6+set_id*16+12], codeword_reg14[256*6+set_id*16+12], codeword_reg13[256*6+set_id*16+12], codeword_reg12[256*6+set_id*16+12], codeword_reg11[256*6+set_id*16+12], codeword_reg10[256*6+set_id*16+12], codeword_reg9[256*6+set_id*16+12], codeword_reg8[256*6+set_id*16+12], codeword_reg7[256*6+set_id*16+12], codeword_reg6[256*6+set_id*16+12], codeword_reg5[256*6+set_id*16+12], codeword_reg4[256*6+set_id*16+12], codeword_reg3[256*6+set_id*16+12], codeword_reg2[256*6+set_id*16+12], codeword_reg1[256*6+set_id*16+12], codeword_reg16[256*5+set_id*16+12], codeword_reg15[256*5+set_id*16+12], codeword_reg14[256*5+set_id*16+12], codeword_reg13[256*5+set_id*16+12], codeword_reg12[256*5+set_id*16+12], codeword_reg11[256*5+set_id*16+12], codeword_reg10[256*5+set_id*16+12], codeword_reg9[256*5+set_id*16+12], codeword_reg8[256*5+set_id*16+12], codeword_reg7[256*5+set_id*16+12], codeword_reg6[256*5+set_id*16+12], codeword_reg5[256*5+set_id*16+12], codeword_reg4[256*5+set_id*16+12], codeword_reg3[256*5+set_id*16+12], codeword_reg2[256*5+set_id*16+12], codeword_reg1[256*5+set_id*16+12], codeword_reg16[256*4+set_id*16+12], codeword_reg15[256*4+set_id*16+12], codeword_reg14[256*4+set_id*16+12], codeword_reg13[256*4+set_id*16+12], codeword_reg12[256*4+set_id*16+12], codeword_reg11[256*4+set_id*16+12], codeword_reg10[256*4+set_id*16+12], codeword_reg9[256*4+set_id*16+12], codeword_reg8[256*4+set_id*16+12], codeword_reg7[256*4+set_id*16+12], codeword_reg6[256*4+set_id*16+12], codeword_reg5[256*4+set_id*16+12], codeword_reg4[256*4+set_id*16+12], codeword_reg3[256*4+set_id*16+12], codeword_reg2[256*4+set_id*16+12], codeword_reg1[256*4+set_id*16+12], codeword_reg16[256*3+set_id*16+12], codeword_reg15[256*3+set_id*16+12], codeword_reg14[256*3+set_id*16+12], codeword_reg13[256*3+set_id*16+12], codeword_reg12[256*3+set_id*16+12], codeword_reg11[256*3+set_id*16+12], codeword_reg10[256*3+set_id*16+12], codeword_reg9[256*3+set_id*16+12], codeword_reg8[256*3+set_id*16+12], codeword_reg7[256*3+set_id*16+12], codeword_reg6[256*3+set_id*16+12], codeword_reg5[256*3+set_id*16+12], codeword_reg4[256*3+set_id*16+12], codeword_reg3[256*3+set_id*16+12], codeword_reg2[256*3+set_id*16+12], codeword_reg1[256*3+set_id*16+12], codeword_reg16[256*2+set_id*16+12], codeword_reg15[256*2+set_id*16+12], codeword_reg14[256*2+set_id*16+12], codeword_reg13[256*2+set_id*16+12], codeword_reg12[256*2+set_id*16+12], codeword_reg11[256*2+set_id*16+12], codeword_reg10[256*2+set_id*16+12], codeword_reg9[256*2+set_id*16+12], codeword_reg8[256*2+set_id*16+12], codeword_reg7[256*2+set_id*16+12], codeword_reg6[256*2+set_id*16+12], codeword_reg5[256*2+set_id*16+12], codeword_reg4[256*2+set_id*16+12], codeword_reg3[256*2+set_id*16+12], codeword_reg2[256*2+set_id*16+12], codeword_reg1[256*2+set_id*16+12], codeword_reg16[256*1+set_id*16+12], codeword_reg15[256*1+set_id*16+12], codeword_reg14[256*1+set_id*16+12], codeword_reg13[256*1+set_id*16+12], codeword_reg12[256*1+set_id*16+12], codeword_reg11[256*1+set_id*16+12], codeword_reg10[256*1+set_id*16+12], codeword_reg9[256*1+set_id*16+12], codeword_reg8[256*1+set_id*16+12], codeword_reg7[256*1+set_id*16+12], codeword_reg6[256*1+set_id*16+12], codeword_reg5[256*1+set_id*16+12], codeword_reg4[256*1+set_id*16+12], codeword_reg3[256*1+set_id*16+12], codeword_reg2[256*1+set_id*16+12], codeword_reg1[256*1+set_id*16+12], codeword_reg16[256*0+set_id*16+12], codeword_reg15[256*0+set_id*16+12], codeword_reg14[256*0+set_id*16+12], codeword_reg13[256*0+set_id*16+12], codeword_reg12[256*0+set_id*16+12], codeword_reg11[256*0+set_id*16+12], codeword_reg10[256*0+set_id*16+12], codeword_reg9[256*0+set_id*16+12], codeword_reg8[256*0+set_id*16+12], codeword_reg7[256*0+set_id*16+12], codeword_reg6[256*0+set_id*16+12], codeword_reg5[256*0+set_id*16+12], codeword_reg4[256*0+set_id*16+12], codeword_reg3[256*0+set_id*16+12], codeword_reg2[256*0+set_id*16+12], codeword_reg1[256*0+set_id*16+12]};
                            in_bits14 <= {codeword_reg16[256*14+set_id*16+13], codeword_reg15[256*14+set_id*16+13], codeword_reg14[256*14+set_id*16+13], codeword_reg13[256*14+set_id*16+13], codeword_reg12[256*14+set_id*16+13], codeword_reg11[256*14+set_id*16+13], codeword_reg10[256*14+set_id*16+13], codeword_reg9[256*14+set_id*16+13], codeword_reg8[256*14+set_id*16+13], codeword_reg7[256*14+set_id*16+13], codeword_reg6[256*14+set_id*16+13], codeword_reg5[256*14+set_id*16+13], codeword_reg4[256*14+set_id*16+13], codeword_reg3[256*14+set_id*16+13], codeword_reg2[256*14+set_id*16+13], codeword_reg1[256*14+set_id*16+13], codeword_reg16[256*13+set_id*16+13], codeword_reg15[256*13+set_id*16+13], codeword_reg14[256*13+set_id*16+13], codeword_reg13[256*13+set_id*16+13], codeword_reg12[256*13+set_id*16+13], codeword_reg11[256*13+set_id*16+13], codeword_reg10[256*13+set_id*16+13], codeword_reg9[256*13+set_id*16+13], codeword_reg8[256*13+set_id*16+13], codeword_reg7[256*13+set_id*16+13], codeword_reg6[256*13+set_id*16+13], codeword_reg5[256*13+set_id*16+13], codeword_reg4[256*13+set_id*16+13], codeword_reg3[256*13+set_id*16+13], codeword_reg2[256*13+set_id*16+13], codeword_reg1[256*13+set_id*16+13], codeword_reg16[256*12+set_id*16+13], codeword_reg15[256*12+set_id*16+13], codeword_reg14[256*12+set_id*16+13], codeword_reg13[256*12+set_id*16+13], codeword_reg12[256*12+set_id*16+13], codeword_reg11[256*12+set_id*16+13], codeword_reg10[256*12+set_id*16+13], codeword_reg9[256*12+set_id*16+13], codeword_reg8[256*12+set_id*16+13], codeword_reg7[256*12+set_id*16+13], codeword_reg6[256*12+set_id*16+13], codeword_reg5[256*12+set_id*16+13], codeword_reg4[256*12+set_id*16+13], codeword_reg3[256*12+set_id*16+13], codeword_reg2[256*12+set_id*16+13], codeword_reg1[256*12+set_id*16+13], codeword_reg16[256*11+set_id*16+13], codeword_reg15[256*11+set_id*16+13], codeword_reg14[256*11+set_id*16+13], codeword_reg13[256*11+set_id*16+13], codeword_reg12[256*11+set_id*16+13], codeword_reg11[256*11+set_id*16+13], codeword_reg10[256*11+set_id*16+13], codeword_reg9[256*11+set_id*16+13], codeword_reg8[256*11+set_id*16+13], codeword_reg7[256*11+set_id*16+13], codeword_reg6[256*11+set_id*16+13], codeword_reg5[256*11+set_id*16+13], codeword_reg4[256*11+set_id*16+13], codeword_reg3[256*11+set_id*16+13], codeword_reg2[256*11+set_id*16+13], codeword_reg1[256*11+set_id*16+13], codeword_reg16[256*10+set_id*16+13], codeword_reg15[256*10+set_id*16+13], codeword_reg14[256*10+set_id*16+13], codeword_reg13[256*10+set_id*16+13], codeword_reg12[256*10+set_id*16+13], codeword_reg11[256*10+set_id*16+13], codeword_reg10[256*10+set_id*16+13], codeword_reg9[256*10+set_id*16+13], codeword_reg8[256*10+set_id*16+13], codeword_reg7[256*10+set_id*16+13], codeword_reg6[256*10+set_id*16+13], codeword_reg5[256*10+set_id*16+13], codeword_reg4[256*10+set_id*16+13], codeword_reg3[256*10+set_id*16+13], codeword_reg2[256*10+set_id*16+13], codeword_reg1[256*10+set_id*16+13], codeword_reg16[256*9+set_id*16+13], codeword_reg15[256*9+set_id*16+13], codeword_reg14[256*9+set_id*16+13], codeword_reg13[256*9+set_id*16+13], codeword_reg12[256*9+set_id*16+13], codeword_reg11[256*9+set_id*16+13], codeword_reg10[256*9+set_id*16+13], codeword_reg9[256*9+set_id*16+13], codeword_reg8[256*9+set_id*16+13], codeword_reg7[256*9+set_id*16+13], codeword_reg6[256*9+set_id*16+13], codeword_reg5[256*9+set_id*16+13], codeword_reg4[256*9+set_id*16+13], codeword_reg3[256*9+set_id*16+13], codeword_reg2[256*9+set_id*16+13], codeword_reg1[256*9+set_id*16+13], codeword_reg16[256*8+set_id*16+13], codeword_reg15[256*8+set_id*16+13], codeword_reg14[256*8+set_id*16+13], codeword_reg13[256*8+set_id*16+13], codeword_reg12[256*8+set_id*16+13], codeword_reg11[256*8+set_id*16+13], codeword_reg10[256*8+set_id*16+13], codeword_reg9[256*8+set_id*16+13], codeword_reg8[256*8+set_id*16+13], codeword_reg7[256*8+set_id*16+13], codeword_reg6[256*8+set_id*16+13], codeword_reg5[256*8+set_id*16+13], codeword_reg4[256*8+set_id*16+13], codeword_reg3[256*8+set_id*16+13], codeword_reg2[256*8+set_id*16+13], codeword_reg1[256*8+set_id*16+13], codeword_reg16[256*7+set_id*16+13], codeword_reg15[256*7+set_id*16+13], codeword_reg14[256*7+set_id*16+13], codeword_reg13[256*7+set_id*16+13], codeword_reg12[256*7+set_id*16+13], codeword_reg11[256*7+set_id*16+13], codeword_reg10[256*7+set_id*16+13], codeword_reg9[256*7+set_id*16+13], codeword_reg8[256*7+set_id*16+13], codeword_reg7[256*7+set_id*16+13], codeword_reg6[256*7+set_id*16+13], codeword_reg5[256*7+set_id*16+13], codeword_reg4[256*7+set_id*16+13], codeword_reg3[256*7+set_id*16+13], codeword_reg2[256*7+set_id*16+13], codeword_reg1[256*7+set_id*16+13], codeword_reg16[256*6+set_id*16+13], codeword_reg15[256*6+set_id*16+13], codeword_reg14[256*6+set_id*16+13], codeword_reg13[256*6+set_id*16+13], codeword_reg12[256*6+set_id*16+13], codeword_reg11[256*6+set_id*16+13], codeword_reg10[256*6+set_id*16+13], codeword_reg9[256*6+set_id*16+13], codeword_reg8[256*6+set_id*16+13], codeword_reg7[256*6+set_id*16+13], codeword_reg6[256*6+set_id*16+13], codeword_reg5[256*6+set_id*16+13], codeword_reg4[256*6+set_id*16+13], codeword_reg3[256*6+set_id*16+13], codeword_reg2[256*6+set_id*16+13], codeword_reg1[256*6+set_id*16+13], codeword_reg16[256*5+set_id*16+13], codeword_reg15[256*5+set_id*16+13], codeword_reg14[256*5+set_id*16+13], codeword_reg13[256*5+set_id*16+13], codeword_reg12[256*5+set_id*16+13], codeword_reg11[256*5+set_id*16+13], codeword_reg10[256*5+set_id*16+13], codeword_reg9[256*5+set_id*16+13], codeword_reg8[256*5+set_id*16+13], codeword_reg7[256*5+set_id*16+13], codeword_reg6[256*5+set_id*16+13], codeword_reg5[256*5+set_id*16+13], codeword_reg4[256*5+set_id*16+13], codeword_reg3[256*5+set_id*16+13], codeword_reg2[256*5+set_id*16+13], codeword_reg1[256*5+set_id*16+13], codeword_reg16[256*4+set_id*16+13], codeword_reg15[256*4+set_id*16+13], codeword_reg14[256*4+set_id*16+13], codeword_reg13[256*4+set_id*16+13], codeword_reg12[256*4+set_id*16+13], codeword_reg11[256*4+set_id*16+13], codeword_reg10[256*4+set_id*16+13], codeword_reg9[256*4+set_id*16+13], codeword_reg8[256*4+set_id*16+13], codeword_reg7[256*4+set_id*16+13], codeword_reg6[256*4+set_id*16+13], codeword_reg5[256*4+set_id*16+13], codeword_reg4[256*4+set_id*16+13], codeword_reg3[256*4+set_id*16+13], codeword_reg2[256*4+set_id*16+13], codeword_reg1[256*4+set_id*16+13], codeword_reg16[256*3+set_id*16+13], codeword_reg15[256*3+set_id*16+13], codeword_reg14[256*3+set_id*16+13], codeword_reg13[256*3+set_id*16+13], codeword_reg12[256*3+set_id*16+13], codeword_reg11[256*3+set_id*16+13], codeword_reg10[256*3+set_id*16+13], codeword_reg9[256*3+set_id*16+13], codeword_reg8[256*3+set_id*16+13], codeword_reg7[256*3+set_id*16+13], codeword_reg6[256*3+set_id*16+13], codeword_reg5[256*3+set_id*16+13], codeword_reg4[256*3+set_id*16+13], codeword_reg3[256*3+set_id*16+13], codeword_reg2[256*3+set_id*16+13], codeword_reg1[256*3+set_id*16+13], codeword_reg16[256*2+set_id*16+13], codeword_reg15[256*2+set_id*16+13], codeword_reg14[256*2+set_id*16+13], codeword_reg13[256*2+set_id*16+13], codeword_reg12[256*2+set_id*16+13], codeword_reg11[256*2+set_id*16+13], codeword_reg10[256*2+set_id*16+13], codeword_reg9[256*2+set_id*16+13], codeword_reg8[256*2+set_id*16+13], codeword_reg7[256*2+set_id*16+13], codeword_reg6[256*2+set_id*16+13], codeword_reg5[256*2+set_id*16+13], codeword_reg4[256*2+set_id*16+13], codeword_reg3[256*2+set_id*16+13], codeword_reg2[256*2+set_id*16+13], codeword_reg1[256*2+set_id*16+13], codeword_reg16[256*1+set_id*16+13], codeword_reg15[256*1+set_id*16+13], codeword_reg14[256*1+set_id*16+13], codeword_reg13[256*1+set_id*16+13], codeword_reg12[256*1+set_id*16+13], codeword_reg11[256*1+set_id*16+13], codeword_reg10[256*1+set_id*16+13], codeword_reg9[256*1+set_id*16+13], codeword_reg8[256*1+set_id*16+13], codeword_reg7[256*1+set_id*16+13], codeword_reg6[256*1+set_id*16+13], codeword_reg5[256*1+set_id*16+13], codeword_reg4[256*1+set_id*16+13], codeword_reg3[256*1+set_id*16+13], codeword_reg2[256*1+set_id*16+13], codeword_reg1[256*1+set_id*16+13], codeword_reg16[256*0+set_id*16+13], codeword_reg15[256*0+set_id*16+13], codeword_reg14[256*0+set_id*16+13], codeword_reg13[256*0+set_id*16+13], codeword_reg12[256*0+set_id*16+13], codeword_reg11[256*0+set_id*16+13], codeword_reg10[256*0+set_id*16+13], codeword_reg9[256*0+set_id*16+13], codeword_reg8[256*0+set_id*16+13], codeword_reg7[256*0+set_id*16+13], codeword_reg6[256*0+set_id*16+13], codeword_reg5[256*0+set_id*16+13], codeword_reg4[256*0+set_id*16+13], codeword_reg3[256*0+set_id*16+13], codeword_reg2[256*0+set_id*16+13], codeword_reg1[256*0+set_id*16+13]};
                            in_bits15 <= {codeword_reg16[256*14+set_id*16+14], codeword_reg15[256*14+set_id*16+14], codeword_reg14[256*14+set_id*16+14], codeword_reg13[256*14+set_id*16+14], codeword_reg12[256*14+set_id*16+14], codeword_reg11[256*14+set_id*16+14], codeword_reg10[256*14+set_id*16+14], codeword_reg9[256*14+set_id*16+14], codeword_reg8[256*14+set_id*16+14], codeword_reg7[256*14+set_id*16+14], codeword_reg6[256*14+set_id*16+14], codeword_reg5[256*14+set_id*16+14], codeword_reg4[256*14+set_id*16+14], codeword_reg3[256*14+set_id*16+14], codeword_reg2[256*14+set_id*16+14], codeword_reg1[256*14+set_id*16+14], codeword_reg16[256*13+set_id*16+14], codeword_reg15[256*13+set_id*16+14], codeword_reg14[256*13+set_id*16+14], codeword_reg13[256*13+set_id*16+14], codeword_reg12[256*13+set_id*16+14], codeword_reg11[256*13+set_id*16+14], codeword_reg10[256*13+set_id*16+14], codeword_reg9[256*13+set_id*16+14], codeword_reg8[256*13+set_id*16+14], codeword_reg7[256*13+set_id*16+14], codeword_reg6[256*13+set_id*16+14], codeword_reg5[256*13+set_id*16+14], codeword_reg4[256*13+set_id*16+14], codeword_reg3[256*13+set_id*16+14], codeword_reg2[256*13+set_id*16+14], codeword_reg1[256*13+set_id*16+14], codeword_reg16[256*12+set_id*16+14], codeword_reg15[256*12+set_id*16+14], codeword_reg14[256*12+set_id*16+14], codeword_reg13[256*12+set_id*16+14], codeword_reg12[256*12+set_id*16+14], codeword_reg11[256*12+set_id*16+14], codeword_reg10[256*12+set_id*16+14], codeword_reg9[256*12+set_id*16+14], codeword_reg8[256*12+set_id*16+14], codeword_reg7[256*12+set_id*16+14], codeword_reg6[256*12+set_id*16+14], codeword_reg5[256*12+set_id*16+14], codeword_reg4[256*12+set_id*16+14], codeword_reg3[256*12+set_id*16+14], codeword_reg2[256*12+set_id*16+14], codeword_reg1[256*12+set_id*16+14], codeword_reg16[256*11+set_id*16+14], codeword_reg15[256*11+set_id*16+14], codeword_reg14[256*11+set_id*16+14], codeword_reg13[256*11+set_id*16+14], codeword_reg12[256*11+set_id*16+14], codeword_reg11[256*11+set_id*16+14], codeword_reg10[256*11+set_id*16+14], codeword_reg9[256*11+set_id*16+14], codeword_reg8[256*11+set_id*16+14], codeword_reg7[256*11+set_id*16+14], codeword_reg6[256*11+set_id*16+14], codeword_reg5[256*11+set_id*16+14], codeword_reg4[256*11+set_id*16+14], codeword_reg3[256*11+set_id*16+14], codeword_reg2[256*11+set_id*16+14], codeword_reg1[256*11+set_id*16+14], codeword_reg16[256*10+set_id*16+14], codeword_reg15[256*10+set_id*16+14], codeword_reg14[256*10+set_id*16+14], codeword_reg13[256*10+set_id*16+14], codeword_reg12[256*10+set_id*16+14], codeword_reg11[256*10+set_id*16+14], codeword_reg10[256*10+set_id*16+14], codeword_reg9[256*10+set_id*16+14], codeword_reg8[256*10+set_id*16+14], codeword_reg7[256*10+set_id*16+14], codeword_reg6[256*10+set_id*16+14], codeword_reg5[256*10+set_id*16+14], codeword_reg4[256*10+set_id*16+14], codeword_reg3[256*10+set_id*16+14], codeword_reg2[256*10+set_id*16+14], codeword_reg1[256*10+set_id*16+14], codeword_reg16[256*9+set_id*16+14], codeword_reg15[256*9+set_id*16+14], codeword_reg14[256*9+set_id*16+14], codeword_reg13[256*9+set_id*16+14], codeword_reg12[256*9+set_id*16+14], codeword_reg11[256*9+set_id*16+14], codeword_reg10[256*9+set_id*16+14], codeword_reg9[256*9+set_id*16+14], codeword_reg8[256*9+set_id*16+14], codeword_reg7[256*9+set_id*16+14], codeword_reg6[256*9+set_id*16+14], codeword_reg5[256*9+set_id*16+14], codeword_reg4[256*9+set_id*16+14], codeword_reg3[256*9+set_id*16+14], codeword_reg2[256*9+set_id*16+14], codeword_reg1[256*9+set_id*16+14], codeword_reg16[256*8+set_id*16+14], codeword_reg15[256*8+set_id*16+14], codeword_reg14[256*8+set_id*16+14], codeword_reg13[256*8+set_id*16+14], codeword_reg12[256*8+set_id*16+14], codeword_reg11[256*8+set_id*16+14], codeword_reg10[256*8+set_id*16+14], codeword_reg9[256*8+set_id*16+14], codeword_reg8[256*8+set_id*16+14], codeword_reg7[256*8+set_id*16+14], codeword_reg6[256*8+set_id*16+14], codeword_reg5[256*8+set_id*16+14], codeword_reg4[256*8+set_id*16+14], codeword_reg3[256*8+set_id*16+14], codeword_reg2[256*8+set_id*16+14], codeword_reg1[256*8+set_id*16+14], codeword_reg16[256*7+set_id*16+14], codeword_reg15[256*7+set_id*16+14], codeword_reg14[256*7+set_id*16+14], codeword_reg13[256*7+set_id*16+14], codeword_reg12[256*7+set_id*16+14], codeword_reg11[256*7+set_id*16+14], codeword_reg10[256*7+set_id*16+14], codeword_reg9[256*7+set_id*16+14], codeword_reg8[256*7+set_id*16+14], codeword_reg7[256*7+set_id*16+14], codeword_reg6[256*7+set_id*16+14], codeword_reg5[256*7+set_id*16+14], codeword_reg4[256*7+set_id*16+14], codeword_reg3[256*7+set_id*16+14], codeword_reg2[256*7+set_id*16+14], codeword_reg1[256*7+set_id*16+14], codeword_reg16[256*6+set_id*16+14], codeword_reg15[256*6+set_id*16+14], codeword_reg14[256*6+set_id*16+14], codeword_reg13[256*6+set_id*16+14], codeword_reg12[256*6+set_id*16+14], codeword_reg11[256*6+set_id*16+14], codeword_reg10[256*6+set_id*16+14], codeword_reg9[256*6+set_id*16+14], codeword_reg8[256*6+set_id*16+14], codeword_reg7[256*6+set_id*16+14], codeword_reg6[256*6+set_id*16+14], codeword_reg5[256*6+set_id*16+14], codeword_reg4[256*6+set_id*16+14], codeword_reg3[256*6+set_id*16+14], codeword_reg2[256*6+set_id*16+14], codeword_reg1[256*6+set_id*16+14], codeword_reg16[256*5+set_id*16+14], codeword_reg15[256*5+set_id*16+14], codeword_reg14[256*5+set_id*16+14], codeword_reg13[256*5+set_id*16+14], codeword_reg12[256*5+set_id*16+14], codeword_reg11[256*5+set_id*16+14], codeword_reg10[256*5+set_id*16+14], codeword_reg9[256*5+set_id*16+14], codeword_reg8[256*5+set_id*16+14], codeword_reg7[256*5+set_id*16+14], codeword_reg6[256*5+set_id*16+14], codeword_reg5[256*5+set_id*16+14], codeword_reg4[256*5+set_id*16+14], codeword_reg3[256*5+set_id*16+14], codeword_reg2[256*5+set_id*16+14], codeword_reg1[256*5+set_id*16+14], codeword_reg16[256*4+set_id*16+14], codeword_reg15[256*4+set_id*16+14], codeword_reg14[256*4+set_id*16+14], codeword_reg13[256*4+set_id*16+14], codeword_reg12[256*4+set_id*16+14], codeword_reg11[256*4+set_id*16+14], codeword_reg10[256*4+set_id*16+14], codeword_reg9[256*4+set_id*16+14], codeword_reg8[256*4+set_id*16+14], codeword_reg7[256*4+set_id*16+14], codeword_reg6[256*4+set_id*16+14], codeword_reg5[256*4+set_id*16+14], codeword_reg4[256*4+set_id*16+14], codeword_reg3[256*4+set_id*16+14], codeword_reg2[256*4+set_id*16+14], codeword_reg1[256*4+set_id*16+14], codeword_reg16[256*3+set_id*16+14], codeword_reg15[256*3+set_id*16+14], codeword_reg14[256*3+set_id*16+14], codeword_reg13[256*3+set_id*16+14], codeword_reg12[256*3+set_id*16+14], codeword_reg11[256*3+set_id*16+14], codeword_reg10[256*3+set_id*16+14], codeword_reg9[256*3+set_id*16+14], codeword_reg8[256*3+set_id*16+14], codeword_reg7[256*3+set_id*16+14], codeword_reg6[256*3+set_id*16+14], codeword_reg5[256*3+set_id*16+14], codeword_reg4[256*3+set_id*16+14], codeword_reg3[256*3+set_id*16+14], codeword_reg2[256*3+set_id*16+14], codeword_reg1[256*3+set_id*16+14], codeword_reg16[256*2+set_id*16+14], codeword_reg15[256*2+set_id*16+14], codeword_reg14[256*2+set_id*16+14], codeword_reg13[256*2+set_id*16+14], codeword_reg12[256*2+set_id*16+14], codeword_reg11[256*2+set_id*16+14], codeword_reg10[256*2+set_id*16+14], codeword_reg9[256*2+set_id*16+14], codeword_reg8[256*2+set_id*16+14], codeword_reg7[256*2+set_id*16+14], codeword_reg6[256*2+set_id*16+14], codeword_reg5[256*2+set_id*16+14], codeword_reg4[256*2+set_id*16+14], codeword_reg3[256*2+set_id*16+14], codeword_reg2[256*2+set_id*16+14], codeword_reg1[256*2+set_id*16+14], codeword_reg16[256*1+set_id*16+14], codeword_reg15[256*1+set_id*16+14], codeword_reg14[256*1+set_id*16+14], codeword_reg13[256*1+set_id*16+14], codeword_reg12[256*1+set_id*16+14], codeword_reg11[256*1+set_id*16+14], codeword_reg10[256*1+set_id*16+14], codeword_reg9[256*1+set_id*16+14], codeword_reg8[256*1+set_id*16+14], codeword_reg7[256*1+set_id*16+14], codeword_reg6[256*1+set_id*16+14], codeword_reg5[256*1+set_id*16+14], codeword_reg4[256*1+set_id*16+14], codeword_reg3[256*1+set_id*16+14], codeword_reg2[256*1+set_id*16+14], codeword_reg1[256*1+set_id*16+14], codeword_reg16[256*0+set_id*16+14], codeword_reg15[256*0+set_id*16+14], codeword_reg14[256*0+set_id*16+14], codeword_reg13[256*0+set_id*16+14], codeword_reg12[256*0+set_id*16+14], codeword_reg11[256*0+set_id*16+14], codeword_reg10[256*0+set_id*16+14], codeword_reg9[256*0+set_id*16+14], codeword_reg8[256*0+set_id*16+14], codeword_reg7[256*0+set_id*16+14], codeword_reg6[256*0+set_id*16+14], codeword_reg5[256*0+set_id*16+14], codeword_reg4[256*0+set_id*16+14], codeword_reg3[256*0+set_id*16+14], codeword_reg2[256*0+set_id*16+14], codeword_reg1[256*0+set_id*16+14]};
                            in_bits16 <= {codeword_reg16[256*14+set_id*16+15], codeword_reg15[256*14+set_id*16+15], codeword_reg14[256*14+set_id*16+15], codeword_reg13[256*14+set_id*16+15], codeword_reg12[256*14+set_id*16+15], codeword_reg11[256*14+set_id*16+15], codeword_reg10[256*14+set_id*16+15], codeword_reg9[256*14+set_id*16+15], codeword_reg8[256*14+set_id*16+15], codeword_reg7[256*14+set_id*16+15], codeword_reg6[256*14+set_id*16+15], codeword_reg5[256*14+set_id*16+15], codeword_reg4[256*14+set_id*16+15], codeword_reg3[256*14+set_id*16+15], codeword_reg2[256*14+set_id*16+15], codeword_reg1[256*14+set_id*16+15], codeword_reg16[256*13+set_id*16+15], codeword_reg15[256*13+set_id*16+15], codeword_reg14[256*13+set_id*16+15], codeword_reg13[256*13+set_id*16+15], codeword_reg12[256*13+set_id*16+15], codeword_reg11[256*13+set_id*16+15], codeword_reg10[256*13+set_id*16+15], codeword_reg9[256*13+set_id*16+15], codeword_reg8[256*13+set_id*16+15], codeword_reg7[256*13+set_id*16+15], codeword_reg6[256*13+set_id*16+15], codeword_reg5[256*13+set_id*16+15], codeword_reg4[256*13+set_id*16+15], codeword_reg3[256*13+set_id*16+15], codeword_reg2[256*13+set_id*16+15], codeword_reg1[256*13+set_id*16+15], codeword_reg16[256*12+set_id*16+15], codeword_reg15[256*12+set_id*16+15], codeword_reg14[256*12+set_id*16+15], codeword_reg13[256*12+set_id*16+15], codeword_reg12[256*12+set_id*16+15], codeword_reg11[256*12+set_id*16+15], codeword_reg10[256*12+set_id*16+15], codeword_reg9[256*12+set_id*16+15], codeword_reg8[256*12+set_id*16+15], codeword_reg7[256*12+set_id*16+15], codeword_reg6[256*12+set_id*16+15], codeword_reg5[256*12+set_id*16+15], codeword_reg4[256*12+set_id*16+15], codeword_reg3[256*12+set_id*16+15], codeword_reg2[256*12+set_id*16+15], codeword_reg1[256*12+set_id*16+15], codeword_reg16[256*11+set_id*16+15], codeword_reg15[256*11+set_id*16+15], codeword_reg14[256*11+set_id*16+15], codeword_reg13[256*11+set_id*16+15], codeword_reg12[256*11+set_id*16+15], codeword_reg11[256*11+set_id*16+15], codeword_reg10[256*11+set_id*16+15], codeword_reg9[256*11+set_id*16+15], codeword_reg8[256*11+set_id*16+15], codeword_reg7[256*11+set_id*16+15], codeword_reg6[256*11+set_id*16+15], codeword_reg5[256*11+set_id*16+15], codeword_reg4[256*11+set_id*16+15], codeword_reg3[256*11+set_id*16+15], codeword_reg2[256*11+set_id*16+15], codeword_reg1[256*11+set_id*16+15], codeword_reg16[256*10+set_id*16+15], codeword_reg15[256*10+set_id*16+15], codeword_reg14[256*10+set_id*16+15], codeword_reg13[256*10+set_id*16+15], codeword_reg12[256*10+set_id*16+15], codeword_reg11[256*10+set_id*16+15], codeword_reg10[256*10+set_id*16+15], codeword_reg9[256*10+set_id*16+15], codeword_reg8[256*10+set_id*16+15], codeword_reg7[256*10+set_id*16+15], codeword_reg6[256*10+set_id*16+15], codeword_reg5[256*10+set_id*16+15], codeword_reg4[256*10+set_id*16+15], codeword_reg3[256*10+set_id*16+15], codeword_reg2[256*10+set_id*16+15], codeword_reg1[256*10+set_id*16+15], codeword_reg16[256*9+set_id*16+15], codeword_reg15[256*9+set_id*16+15], codeword_reg14[256*9+set_id*16+15], codeword_reg13[256*9+set_id*16+15], codeword_reg12[256*9+set_id*16+15], codeword_reg11[256*9+set_id*16+15], codeword_reg10[256*9+set_id*16+15], codeword_reg9[256*9+set_id*16+15], codeword_reg8[256*9+set_id*16+15], codeword_reg7[256*9+set_id*16+15], codeword_reg6[256*9+set_id*16+15], codeword_reg5[256*9+set_id*16+15], codeword_reg4[256*9+set_id*16+15], codeword_reg3[256*9+set_id*16+15], codeword_reg2[256*9+set_id*16+15], codeword_reg1[256*9+set_id*16+15], codeword_reg16[256*8+set_id*16+15], codeword_reg15[256*8+set_id*16+15], codeword_reg14[256*8+set_id*16+15], codeword_reg13[256*8+set_id*16+15], codeword_reg12[256*8+set_id*16+15], codeword_reg11[256*8+set_id*16+15], codeword_reg10[256*8+set_id*16+15], codeword_reg9[256*8+set_id*16+15], codeword_reg8[256*8+set_id*16+15], codeword_reg7[256*8+set_id*16+15], codeword_reg6[256*8+set_id*16+15], codeword_reg5[256*8+set_id*16+15], codeword_reg4[256*8+set_id*16+15], codeword_reg3[256*8+set_id*16+15], codeword_reg2[256*8+set_id*16+15], codeword_reg1[256*8+set_id*16+15], codeword_reg16[256*7+set_id*16+15], codeword_reg15[256*7+set_id*16+15], codeword_reg14[256*7+set_id*16+15], codeword_reg13[256*7+set_id*16+15], codeword_reg12[256*7+set_id*16+15], codeword_reg11[256*7+set_id*16+15], codeword_reg10[256*7+set_id*16+15], codeword_reg9[256*7+set_id*16+15], codeword_reg8[256*7+set_id*16+15], codeword_reg7[256*7+set_id*16+15], codeword_reg6[256*7+set_id*16+15], codeword_reg5[256*7+set_id*16+15], codeword_reg4[256*7+set_id*16+15], codeword_reg3[256*7+set_id*16+15], codeword_reg2[256*7+set_id*16+15], codeword_reg1[256*7+set_id*16+15], codeword_reg16[256*6+set_id*16+15], codeword_reg15[256*6+set_id*16+15], codeword_reg14[256*6+set_id*16+15], codeword_reg13[256*6+set_id*16+15], codeword_reg12[256*6+set_id*16+15], codeword_reg11[256*6+set_id*16+15], codeword_reg10[256*6+set_id*16+15], codeword_reg9[256*6+set_id*16+15], codeword_reg8[256*6+set_id*16+15], codeword_reg7[256*6+set_id*16+15], codeword_reg6[256*6+set_id*16+15], codeword_reg5[256*6+set_id*16+15], codeword_reg4[256*6+set_id*16+15], codeword_reg3[256*6+set_id*16+15], codeword_reg2[256*6+set_id*16+15], codeword_reg1[256*6+set_id*16+15], codeword_reg16[256*5+set_id*16+15], codeword_reg15[256*5+set_id*16+15], codeword_reg14[256*5+set_id*16+15], codeword_reg13[256*5+set_id*16+15], codeword_reg12[256*5+set_id*16+15], codeword_reg11[256*5+set_id*16+15], codeword_reg10[256*5+set_id*16+15], codeword_reg9[256*5+set_id*16+15], codeword_reg8[256*5+set_id*16+15], codeword_reg7[256*5+set_id*16+15], codeword_reg6[256*5+set_id*16+15], codeword_reg5[256*5+set_id*16+15], codeword_reg4[256*5+set_id*16+15], codeword_reg3[256*5+set_id*16+15], codeword_reg2[256*5+set_id*16+15], codeword_reg1[256*5+set_id*16+15], codeword_reg16[256*4+set_id*16+15], codeword_reg15[256*4+set_id*16+15], codeword_reg14[256*4+set_id*16+15], codeword_reg13[256*4+set_id*16+15], codeword_reg12[256*4+set_id*16+15], codeword_reg11[256*4+set_id*16+15], codeword_reg10[256*4+set_id*16+15], codeword_reg9[256*4+set_id*16+15], codeword_reg8[256*4+set_id*16+15], codeword_reg7[256*4+set_id*16+15], codeword_reg6[256*4+set_id*16+15], codeword_reg5[256*4+set_id*16+15], codeword_reg4[256*4+set_id*16+15], codeword_reg3[256*4+set_id*16+15], codeword_reg2[256*4+set_id*16+15], codeword_reg1[256*4+set_id*16+15], codeword_reg16[256*3+set_id*16+15], codeword_reg15[256*3+set_id*16+15], codeword_reg14[256*3+set_id*16+15], codeword_reg13[256*3+set_id*16+15], codeword_reg12[256*3+set_id*16+15], codeword_reg11[256*3+set_id*16+15], codeword_reg10[256*3+set_id*16+15], codeword_reg9[256*3+set_id*16+15], codeword_reg8[256*3+set_id*16+15], codeword_reg7[256*3+set_id*16+15], codeword_reg6[256*3+set_id*16+15], codeword_reg5[256*3+set_id*16+15], codeword_reg4[256*3+set_id*16+15], codeword_reg3[256*3+set_id*16+15], codeword_reg2[256*3+set_id*16+15], codeword_reg1[256*3+set_id*16+15], codeword_reg16[256*2+set_id*16+15], codeword_reg15[256*2+set_id*16+15], codeword_reg14[256*2+set_id*16+15], codeword_reg13[256*2+set_id*16+15], codeword_reg12[256*2+set_id*16+15], codeword_reg11[256*2+set_id*16+15], codeword_reg10[256*2+set_id*16+15], codeword_reg9[256*2+set_id*16+15], codeword_reg8[256*2+set_id*16+15], codeword_reg7[256*2+set_id*16+15], codeword_reg6[256*2+set_id*16+15], codeword_reg5[256*2+set_id*16+15], codeword_reg4[256*2+set_id*16+15], codeword_reg3[256*2+set_id*16+15], codeword_reg2[256*2+set_id*16+15], codeword_reg1[256*2+set_id*16+15], codeword_reg16[256*1+set_id*16+15], codeword_reg15[256*1+set_id*16+15], codeword_reg14[256*1+set_id*16+15], codeword_reg13[256*1+set_id*16+15], codeword_reg12[256*1+set_id*16+15], codeword_reg11[256*1+set_id*16+15], codeword_reg10[256*1+set_id*16+15], codeword_reg9[256*1+set_id*16+15], codeword_reg8[256*1+set_id*16+15], codeword_reg7[256*1+set_id*16+15], codeword_reg6[256*1+set_id*16+15], codeword_reg5[256*1+set_id*16+15], codeword_reg4[256*1+set_id*16+15], codeword_reg3[256*1+set_id*16+15], codeword_reg2[256*1+set_id*16+15], codeword_reg1[256*1+set_id*16+15], codeword_reg16[256*0+set_id*16+15], codeword_reg15[256*0+set_id*16+15], codeword_reg14[256*0+set_id*16+15], codeword_reg13[256*0+set_id*16+15], codeword_reg12[256*0+set_id*16+15], codeword_reg11[256*0+set_id*16+15], codeword_reg10[256*0+set_id*16+15], codeword_reg9[256*0+set_id*16+15], codeword_reg8[256*0+set_id*16+15], codeword_reg7[256*0+set_id*16+15], codeword_reg6[256*0+set_id*16+15], codeword_reg5[256*0+set_id*16+15], codeword_reg4[256*0+set_id*16+15], codeword_reg3[256*0+set_id*16+15], codeword_reg2[256*0+set_id*16+15], codeword_reg1[256*0+set_id*16+15]};
                            
                            // Output the encoded codewords
                            out_codeword1  <= codeword1;
                            out_codeword2  <= codeword2;
                            out_codeword3  <= codeword3;
                            out_codeword4  <= codeword4;
                            out_codeword5  <= codeword5;
                            out_codeword6  <= codeword6;
                            out_codeword7  <= codeword7;
                            out_codeword8  <= codeword8;
                            out_codeword9  <= codeword9;
                            out_codeword10 <= codeword10;
                            out_codeword11 <= codeword11;
                            out_codeword12 <= codeword12;
                            out_codeword13 <= codeword13;
                            out_codeword14 <= codeword14;
                            out_codeword15 <= codeword15;
                            out_codeword16 <= codeword16;
                            
                            // Update the control variables
                            if (col_counter == 5'd1)
                                new1 <= 1'b1;
                            else 
                                new1 <= 1'b0;
                            set_id <= set_id + 4'b1;
                            col_counter <= col_counter + 1;
                            if (col_counter > 5'd0)
                                store <= 1'b1;
                            else
                                store <= 1'b0;
                        
                        // For this range, the input is taken from the bit_gen
                        end else begin
                            
                            // Give generated bits as the input
                            in_bits1  <= bits1;
                            in_bits2  <= bits2;
                            in_bits3  <= bits3;
                            in_bits4  <= bits4;
                            in_bits5  <= bits5;
                            in_bits6  <= bits6;
                            in_bits7  <= bits7;
                            in_bits8  <= bits8;
                            in_bits9  <= bits9;
                            in_bits10 <= bits10;
                            in_bits11 <= bits11;
                            in_bits12 <= bits12;
                            in_bits13 <= bits13;
                            in_bits14 <= bits14;
                            in_bits15 <= bits15;
                            in_bits16 <= bits16;
                            
                            // Output the encoded codewords
                            out_codeword1  <= codeword1;
                            out_codeword2  <= codeword2;
                            out_codeword3  <= codeword3;
                            out_codeword4  <= codeword4;
                            out_codeword5  <= codeword5;
                            out_codeword6  <= codeword6;
                            out_codeword7  <= codeword7;
                            out_codeword8  <= codeword8;
                            out_codeword9  <= codeword9;
                            out_codeword10 <= codeword10;
                            out_codeword11 <= codeword11;
                            out_codeword12 <= codeword12;
                            out_codeword13 <= codeword13;
                            out_codeword14 <= codeword14;
                            out_codeword15 <= codeword15;
                            out_codeword16 <= codeword16;
                            
                            // Update the control variables
                            set_id <= 4'b0;
                            col_counter <= 5'b0;
                            row <= 1'b1;
                            new1 <= 1'b0;
                            store <= 1'b1;
                            start <= 2'b0;
                        end
                    end 
                    //// End of the column encoding ////
                
                // Initiating in_bits
                end else begin 
                    new1 <= 1'b0;
                    
                    in_bits1  <= bits1;
                    in_bits2  <= bits2;
                    in_bits3  <= bits3;
                    in_bits4  <= bits4;
                    in_bits5  <= bits5;
                    in_bits6  <= bits6;
                    in_bits7  <= bits7;
                    in_bits8  <= bits8;
                    in_bits9  <= bits9;
                    in_bits10 <= bits10;
                    in_bits11 <= bits11;
                    in_bits12 <= bits12;
                    in_bits13 <= bits13;
                    in_bits14 <= bits14;
                    in_bits15 <= bits15;
                    in_bits16 <= bits16;
                    
//                    if (start == 2'b0) begin
//                        in_bits1  <= 'bx;
//                        in_bits2  <= 'bx;
//                        in_bits3  <= 'bx;
//                        in_bits4  <= 'bx;
//                        in_bits5  <= 'bx;
//                        in_bits6  <= 'bx;
//                        in_bits7  <= 'bx;
//                        in_bits8  <= 'bx;
//                        in_bits9  <= 'bx;
//                        in_bits10 <= 'bx;
//                        in_bits11 <= 'bx;
//                        in_bits12 <= 'bx;
//                        in_bits13 <= 'bx;
//                        in_bits14 <= 'bx;
//                        in_bits15 <= 'bx;
//                        in_bits16 <= 'bx;
//                    end else begin                
//                        in_bits1  <= bits1;
//                        in_bits2  <= bits2;
//                        in_bits3  <= bits3;
//                        in_bits4  <= bits4;
//                        in_bits5  <= bits5;
//                        in_bits6  <= bits6;
//                        in_bits7  <= bits7;
//                        in_bits8  <= bits8;
//                        in_bits9  <= bits9;
//                        in_bits10 <= bits10;
//                        in_bits11 <= bits11;
//                        in_bits12 <= bits12;
//                        in_bits13 <= bits13;
//                        in_bits14 <= bits14;
//                        in_bits15 <= bits15;
//                        in_bits16 <= bits16;
//                    end
                        
                    new1 <= 1'b0;
                    start <= start + 2'b01;
                    store <= 1'b0;
                end
            //// When the decoding is still in process, the encoding is held
            end else begin // When decoding is still in process
                
                in_bits1  <= 'bx;
                in_bits2  <= 'bx;
                in_bits3  <= 'bx;
                in_bits4  <= 'bx;
                in_bits5  <= 'bx;
                in_bits6  <= 'bx;
                in_bits7  <= 'bx;
                in_bits8  <= 'bx;
                in_bits9  <= 'bx;
                in_bits10 <= 'bx;
                in_bits11 <= 'bx;
                in_bits12 <= 'bx;
                in_bits13 <= 'bx;
                in_bits14 <= 'bx;
                in_bits15 <= 'bx;
                in_bits16 <= 'bx;
            
                out_codeword1  <= 'bx;
                out_codeword2  <= 'bx;
                out_codeword3  <= 'bx;
                out_codeword4  <= 'bx;
                out_codeword5  <= 'bx;
                out_codeword6  <= 'bx;
                out_codeword7  <= 'bx;
                out_codeword8  <= 'bx;
                out_codeword9  <= 'bx;
                out_codeword10 <= 'bx;
                out_codeword11 <= 'bx;
                out_codeword12 <= 'bx;
                out_codeword13 <= 'bx;
                out_codeword14 <= 'bx;
                out_codeword15 <= 'bx;
                out_codeword16 <= 'bx;
                
                new1 <= 1'b0;
                store <= 1'b0;
            end
                
            
        end
    end
endmodule

//always@(posedge clk) begin
//        if (!reset) begin // If reset is 0
//            counter_bit_gen <= 5'b0;
//            counter_hold_bit_gen <= 4'b0;
//            col_id <= 4'b0;
//            start <= 1'b0;
//        end else begin // If reset is 1
//            if (start == 1'b1) begin
//                if (counter_bit_gen < 5'd16) begin // If the bit generation is allowed           
//                    col_id <= col_id + 4'b1;
//                    counter_bit_gen <= counter_bit_gen + 1;
                    
//                    if (counter_bit_gen == 5'd15)
//                        in_bits1  <= bits1;
//                        in_bits2  <= bits2;
//                        in_bits3  <= bits3;
//                        in_bits4  <= bits4;
//                        in_bits5  <= bits5;
//                        in_bits6  <= bits6;
//                        in_bits7  <= bits7;
//                        in_bits8  <= bits8;
//                        in_bits9  <= bits9;
//                        in_bits10 <= bits10;
//                        in_bits11 <= bits11;
//                        in_bits12 <= bits12;
//                        in_bits13 <= bits13;
//                        in_bits14 <= bits14;
//                        in_bits15 <= bits15;
//                        in_bits16 <= bits16;
//                    end else begin
//                        in_bits1  <= bits1;
//                        in_bits2  <= bits2;
//                        in_bits3  <= bits3;
//                        in_bits4  <= bits4;
//                        in_bits5  <= bits5;
//                        in_bits6  <= bits6;
//                        in_bits7  <= bits7;
//                        in_bits8  <= bits8;
//                        in_bits9  <= bits9;
//                        in_bits10 <= bits10;
//                        in_bits11 <= bits11;
//                        in_bits12 <= bits12;
//                        in_bits13 <= bits13;
//                        in_bits14 <= bits14;
//                        in_bits15 <= bits15;
//                        in_bits16 <= bits16;
//                    end
                    
//                    codeword_reg1[(col_id)*n  +: n] <= codeword1;
//                    codeword_reg2[(col_id)*n  +: n] <= codeword2;
//                    codeword_reg3[(col_id)*n  +: n] <= codeword3;
//                    codeword_reg4[(col_id)*n  +: n] <= codeword4;
//                    codeword_reg5[(col_id)*n  +: n] <= codeword5;
//                    codeword_reg6[(col_id)*n  +: n] <= codeword6;
//                    codeword_reg7[(col_id)*n  +: n] <= codeword7;
//                    codeword_reg8[(col_id)*n  +: n] <= codeword8;
//                    codeword_reg9[(col_id)*n  +: n] <= codeword9;
//                    codeword_reg10[(col_id)*n +: n] <= codeword10;
//                    codeword_reg11[(col_id)*n +: n] <= codeword11;
//                    codeword_reg12[(col_id)*n +: n] <= codeword12;
//                    codeword_reg13[(col_id)*n +: n] <= codeword13;
//                    codeword_reg14[(col_id)*n +: n] <= codeword14;
//                    codeword_reg15[(col_id)*n +: n] <= codeword15;
//                    codeword_reg16[(col_id)*n +: n] <= codeword16;
                                   
//                end else begin // If the bit generation is not allowed
//                    if (counter_hold_bit_gen < 4'd15) begin // If the bitgeneration is on hold
//                        counter_hold_bit_gen <= counter_hold_bit_gen + 1;
                        
//                        in_bits1  <= ;
//                        in_bits2  <= ;
//                        in_bits3  <= ;
//                        in_bits4  <= ;
//                        in_bits5  <= ;
//                        in_bits6  <= ;
//                        in_bits7  <= ;
//                        in_bits8  <= ;
//                        in_bits9  <= ;
//                        in_bits10 <= ;
//                        in_bits11 <= ;
//                        in_bits12 <= ;
//                        in_bits13 <= ;
//                        in_bits14 <= ;
//                        in_bits15 <= ;
//                        in_bits16 <= ;
                        
//                    end else begin // If the bit generation is going to be allowed
//                        col_id <= 1'b0;
//                        counter_bit_gen <= 5'b0; 
//                    end    
//                end
//            end else begin
//                in_bits1  <= bits1;
//                in_bits2  <= bits2;
//                in_bits3  <= bits3;
//                in_bits4  <= bits4;
//                in_bits5  <= bits5;
//                in_bits6  <= bits6;
//                in_bits7  <= bits7;
//                in_bits8  <= bits8;
//                in_bits9  <= bits9;
//                in_bits10 <= bits10;
//                in_bits11 <= bits11;
//                in_bits12 <= bits12;
//                in_bits13 <= bits13;
//                in_bits14 <= bits14;
//                in_bits15 <= bits15;
//                in_bits16 <= bits16;
//                counting <= 1'b1;
//            end
//        end
