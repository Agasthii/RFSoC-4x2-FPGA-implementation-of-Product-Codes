`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/11/2024 04:14:15 PM
// Design Name: 
// Module Name: bit_gen_PC
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bit_gen_PC#(
    parameter k = 239
    )(
    input wire clk,
    input wire reset,
    input wire [4095:0] seed,
//     input wire [8191:0] seed,
    output wire [k-1:0] bits1,
    output wire [k-1:0] bits2,
    output wire [k-1:0] bits3,
    output wire [k-1:0] bits4,
    output wire [k-1:0] bits5,
    output wire [k-1:0] bits6,
    output wire [k-1:0] bits7,
    output wire [k-1:0] bits8,
    output wire [k-1:0] bits9,
    output wire [k-1:0] bits10,
    output wire [k-1:0] bits11,
    output wire [k-1:0] bits12,
    output wire [k-1:0] bits13,
    output wire [k-1:0] bits14,
    output wire [k-1:0] bits15,
    output wire [k-1:0] bits16             
    );
    
    // reg [4095:0] lfsr; 
    // reg feedback;

    bit_gen_239 information1(
    .clk(clk),
    .reset(reset),
    .seed(seed[255:0]),
    .bits(bits1)
    );
   bit_gen_239 information2(
    .clk(clk),
    .reset(reset),
    .seed(seed[511:256]),
    .bits(bits2)
    );
   bit_gen_239 information3(
    .clk(clk),
    .reset(reset),
    .seed(seed[767:512]),
    .bits(bits3)
    );
   bit_gen_239 information4(
    .clk(clk),
    .reset(reset),
    .seed(seed[1023:768]),
    .bits(bits4)
    );
   bit_gen_239 information5(
    .clk(clk),
    .reset(reset),
    .seed(seed[1279:1024]),
    .bits(bits5)
    );
   bit_gen_239 information6(
    .clk(clk),
    .reset(reset),
    .seed(seed[1535:1280]),
    .bits(bits6)
    );
   bit_gen_239 information17(
    .clk(clk),
    .reset(reset),
    .seed(seed[1791:1536]),
    .bits(bits7)
    );
   bit_gen_239 information8(
    .clk(clk),
    .reset(reset),
    .seed(seed[2047:1792]),
    .bits(bits8)
    );
   bit_gen_239 information9(
    .clk(clk),
    .reset(reset),
    .seed(seed[2303:2048]),
    .bits(bits9)
    );
   bit_gen_239 information10(
    .clk(clk),
    .reset(reset),
    .seed(seed[2559:2304]),
    .bits(bits10)
    );
   bit_gen_239 information11(
    .clk(clk),
    .reset(reset),
    .seed(seed[2815:2560]),
    .bits(bits11)
    );
   bit_gen_239 information12(
    .clk(clk),
    .reset(reset),
    .seed(seed[3071:2816]),
    .bits(bits12)
    );
   bit_gen_239 information13(
    .clk(clk),
    .reset(reset),
    .seed(seed[3327:3072]),
    .bits(bits13)
    );
   bit_gen_239 information14(
    .clk(clk),
    .reset(reset),
    .seed(seed[3583:3328]),
    .bits(bits14)
    );
   bit_gen_239 information15(
    .clk(clk),
    .reset(reset),
    .seed(seed[3839:3584]),
    .bits(bits15)
    );
   bit_gen_239 information16(
    .clk(clk),
    .reset(reset),
    .seed(seed[4095:3840]),
    .bits(bits16)
    );
    
endmodule


// always @(posedge clk) begin
//         //Update LFSR -> probabilities
//         //Taps at 4096, 4095, 4081, 4069
//         if(reset) begin
//             feedback = lfsr[0];
//             lfsr[4095] = feedback ^ lfsr[4095];
//             lfsr[4094] = feedback ^ lfsr[4094];
//             lfsr[4080] = feedback ^ lfsr[4080];
//             lfsr[4068] = feedback ^ lfsr[4068]; 
//             lfsr = (lfsr >> 1);
//             lfsr[4095] = feedback;
            
//             bits1 <= {lfsr[0], lfsr[1], lfsr[2], lfsr[3], lfsr[4], lfsr[5], lfsr[6], lfsr[7], lfsr[8], lfsr[9], lfsr[10], lfsr[11], lfsr[12], lfsr[13], lfsr[14], lfsr[15], lfsr[16], lfsr[17], lfsr[18], lfsr[19], lfsr[20], lfsr[21], lfsr[22], lfsr[23], lfsr[24], lfsr[25], lfsr[26], lfsr[27], lfsr[28], lfsr[29], lfsr[30], lfsr[31], lfsr[32], lfsr[33], lfsr[34], lfsr[35], lfsr[36], lfsr[37], lfsr[38], lfsr[39], lfsr[40], lfsr[41], lfsr[42], lfsr[43], lfsr[44], lfsr[45], lfsr[46], lfsr[47], lfsr[48], lfsr[49], lfsr[50], lfsr[51], lfsr[52], lfsr[53], lfsr[54], lfsr[55], lfsr[56], lfsr[57], lfsr[58], lfsr[59], lfsr[60], lfsr[61], lfsr[62], lfsr[63], lfsr[64], lfsr[65], lfsr[66], lfsr[67], lfsr[68], lfsr[69], lfsr[70], lfsr[71], lfsr[72], lfsr[73], lfsr[74], lfsr[75], lfsr[76], lfsr[77], lfsr[78], lfsr[79], lfsr[80], lfsr[81], lfsr[82], lfsr[83], lfsr[84], lfsr[85], lfsr[86], lfsr[87], lfsr[88], lfsr[89], lfsr[90], lfsr[91], lfsr[92], lfsr[93], lfsr[94], lfsr[95], lfsr[96], lfsr[97], lfsr[98], lfsr[99], lfsr[100], lfsr[101], lfsr[102], lfsr[103], lfsr[104], lfsr[105], lfsr[106], lfsr[107], lfsr[108], lfsr[109], lfsr[110], lfsr[111], lfsr[112], lfsr[113], lfsr[114], lfsr[115], lfsr[116], lfsr[117], lfsr[118], lfsr[119], lfsr[120], lfsr[121], lfsr[122], lfsr[123], lfsr[124], lfsr[125], lfsr[126], lfsr[127], lfsr[128], lfsr[129], lfsr[130], lfsr[131], lfsr[132], lfsr[133], lfsr[134], lfsr[135], lfsr[136], lfsr[137], lfsr[138], lfsr[139], lfsr[140], lfsr[141], lfsr[142], lfsr[143], lfsr[144], lfsr[145], lfsr[146], lfsr[147], lfsr[148], lfsr[149], lfsr[150], lfsr[151], lfsr[152], lfsr[153], lfsr[154], lfsr[155], lfsr[156], lfsr[157], lfsr[158], lfsr[159], lfsr[160], lfsr[161], lfsr[162], lfsr[163], lfsr[164], lfsr[165], lfsr[166], lfsr[167], lfsr[168], lfsr[169], lfsr[170], lfsr[171], lfsr[172], lfsr[173], lfsr[174], lfsr[175], lfsr[176], lfsr[177], lfsr[178], lfsr[179], lfsr[180], lfsr[181], lfsr[182], lfsr[183], lfsr[184], lfsr[185], lfsr[186], lfsr[187], lfsr[188], lfsr[189], lfsr[190], lfsr[191], lfsr[192], lfsr[193], lfsr[194], lfsr[195], lfsr[196], lfsr[197], lfsr[198], lfsr[199], lfsr[200], lfsr[201], lfsr[202], lfsr[203], lfsr[204], lfsr[205], lfsr[206], lfsr[207], lfsr[208], lfsr[209], lfsr[210], lfsr[211], lfsr[212], lfsr[213], lfsr[214], lfsr[215], lfsr[216], lfsr[217], lfsr[218], lfsr[219], lfsr[220], lfsr[221], lfsr[222], lfsr[223], lfsr[224], lfsr[225], lfsr[226], lfsr[227], lfsr[228], lfsr[229], lfsr[230], lfsr[231], lfsr[232], lfsr[233], lfsr[234], lfsr[235], lfsr[236], lfsr[237], lfsr[238]}; 
//             bits2 <= {lfsr[239], lfsr[240], lfsr[241], lfsr[242], lfsr[243], lfsr[244], lfsr[245], lfsr[246], lfsr[247], lfsr[248], lfsr[249], lfsr[250], lfsr[251], lfsr[252], lfsr[253], lfsr[254], lfsr[255], lfsr[256], lfsr[257], lfsr[258], lfsr[259], lfsr[260], lfsr[261], lfsr[262], lfsr[263], lfsr[264], lfsr[265], lfsr[266], lfsr[267], lfsr[268], lfsr[269], lfsr[270], lfsr[271], lfsr[272], lfsr[273], lfsr[274], lfsr[275], lfsr[276], lfsr[277], lfsr[278], lfsr[279], lfsr[280], lfsr[281], lfsr[282], lfsr[283], lfsr[284], lfsr[285], lfsr[286], lfsr[287], lfsr[288], lfsr[289], lfsr[290], lfsr[291], lfsr[292], lfsr[293], lfsr[294], lfsr[295], lfsr[296], lfsr[297], lfsr[298], lfsr[299], lfsr[300], lfsr[301], lfsr[302], lfsr[303], lfsr[304], lfsr[305], lfsr[306], lfsr[307], lfsr[308], lfsr[309], lfsr[310], lfsr[311], lfsr[312], lfsr[313], lfsr[314], lfsr[315], lfsr[316], lfsr[317], lfsr[318], lfsr[319], lfsr[320], lfsr[321], lfsr[322], lfsr[323], lfsr[324], lfsr[325], lfsr[326], lfsr[327], lfsr[328], lfsr[329], lfsr[330], lfsr[331], lfsr[332], lfsr[333], lfsr[334], lfsr[335], lfsr[336], lfsr[337], lfsr[338], lfsr[339], lfsr[340], lfsr[341], lfsr[342], lfsr[343], lfsr[344], lfsr[345], lfsr[346], lfsr[347], lfsr[348], lfsr[349], lfsr[350], lfsr[351], lfsr[352], lfsr[353], lfsr[354], lfsr[355], lfsr[356], lfsr[357], lfsr[358], lfsr[359], lfsr[360], lfsr[361], lfsr[362], lfsr[363], lfsr[364], lfsr[365], lfsr[366], lfsr[367], lfsr[368], lfsr[369], lfsr[370], lfsr[371], lfsr[372], lfsr[373], lfsr[374], lfsr[375], lfsr[376], lfsr[377], lfsr[378], lfsr[379], lfsr[380], lfsr[381], lfsr[382], lfsr[383], lfsr[384], lfsr[385], lfsr[386], lfsr[387], lfsr[388], lfsr[389], lfsr[390], lfsr[391], lfsr[392], lfsr[393], lfsr[394], lfsr[395], lfsr[396], lfsr[397], lfsr[398], lfsr[399], lfsr[400], lfsr[401], lfsr[402], lfsr[403], lfsr[404], lfsr[405], lfsr[406], lfsr[407], lfsr[408], lfsr[409], lfsr[410], lfsr[411], lfsr[412], lfsr[413], lfsr[414], lfsr[415], lfsr[416], lfsr[417], lfsr[418], lfsr[419], lfsr[420], lfsr[421], lfsr[422], lfsr[423], lfsr[424], lfsr[425], lfsr[426], lfsr[427], lfsr[428], lfsr[429], lfsr[430], lfsr[431], lfsr[432], lfsr[433], lfsr[434], lfsr[435], lfsr[436], lfsr[437], lfsr[438], lfsr[439], lfsr[440], lfsr[441], lfsr[442], lfsr[443], lfsr[444], lfsr[445], lfsr[446], lfsr[447], lfsr[448], lfsr[449], lfsr[450], lfsr[451], lfsr[452], lfsr[453], lfsr[454], lfsr[455], lfsr[456], lfsr[457], lfsr[458], lfsr[459], lfsr[460], lfsr[461], lfsr[462], lfsr[463], lfsr[464], lfsr[465], lfsr[466], lfsr[467], lfsr[468], lfsr[469], lfsr[470], lfsr[471], lfsr[472], lfsr[473], lfsr[474], lfsr[475], lfsr[476], lfsr[477]}; 
//             bits3 <= {lfsr[478], lfsr[479], lfsr[480], lfsr[481], lfsr[482], lfsr[483], lfsr[484], lfsr[485], lfsr[486], lfsr[487], lfsr[488], lfsr[489], lfsr[490], lfsr[491], lfsr[492], lfsr[493], lfsr[494], lfsr[495], lfsr[496], lfsr[497], lfsr[498], lfsr[499], lfsr[500], lfsr[501], lfsr[502], lfsr[503], lfsr[504], lfsr[505], lfsr[506], lfsr[507], lfsr[508], lfsr[509], lfsr[510], lfsr[511], lfsr[512], lfsr[513], lfsr[514], lfsr[515], lfsr[516], lfsr[517], lfsr[518], lfsr[519], lfsr[520], lfsr[521], lfsr[522], lfsr[523], lfsr[524], lfsr[525], lfsr[526], lfsr[527], lfsr[528], lfsr[529], lfsr[530], lfsr[531], lfsr[532], lfsr[533], lfsr[534], lfsr[535], lfsr[536], lfsr[537], lfsr[538], lfsr[539], lfsr[540], lfsr[541], lfsr[542], lfsr[543], lfsr[544], lfsr[545], lfsr[546], lfsr[547], lfsr[548], lfsr[549], lfsr[550], lfsr[551], lfsr[552], lfsr[553], lfsr[554], lfsr[555], lfsr[556], lfsr[557], lfsr[558], lfsr[559], lfsr[560], lfsr[561], lfsr[562], lfsr[563], lfsr[564], lfsr[565], lfsr[566], lfsr[567], lfsr[568], lfsr[569], lfsr[570], lfsr[571], lfsr[572], lfsr[573], lfsr[574], lfsr[575], lfsr[576], lfsr[577], lfsr[578], lfsr[579], lfsr[580], lfsr[581], lfsr[582], lfsr[583], lfsr[584], lfsr[585], lfsr[586], lfsr[587], lfsr[588], lfsr[589], lfsr[590], lfsr[591], lfsr[592], lfsr[593], lfsr[594], lfsr[595], lfsr[596], lfsr[597], lfsr[598], lfsr[599], lfsr[600], lfsr[601], lfsr[602], lfsr[603], lfsr[604], lfsr[605], lfsr[606], lfsr[607], lfsr[608], lfsr[609], lfsr[610], lfsr[611], lfsr[612], lfsr[613], lfsr[614], lfsr[615], lfsr[616], lfsr[617], lfsr[618], lfsr[619], lfsr[620], lfsr[621], lfsr[622], lfsr[623], lfsr[624], lfsr[625], lfsr[626], lfsr[627], lfsr[628], lfsr[629], lfsr[630], lfsr[631], lfsr[632], lfsr[633], lfsr[634], lfsr[635], lfsr[636], lfsr[637], lfsr[638], lfsr[639], lfsr[640], lfsr[641], lfsr[642], lfsr[643], lfsr[644], lfsr[645], lfsr[646], lfsr[647], lfsr[648], lfsr[649], lfsr[650], lfsr[651], lfsr[652], lfsr[653], lfsr[654], lfsr[655], lfsr[656], lfsr[657], lfsr[658], lfsr[659], lfsr[660], lfsr[661], lfsr[662], lfsr[663], lfsr[664], lfsr[665], lfsr[666], lfsr[667], lfsr[668], lfsr[669], lfsr[670], lfsr[671], lfsr[672], lfsr[673], lfsr[674], lfsr[675], lfsr[676], lfsr[677], lfsr[678], lfsr[679], lfsr[680], lfsr[681], lfsr[682], lfsr[683], lfsr[684], lfsr[685], lfsr[686], lfsr[687], lfsr[688], lfsr[689], lfsr[690], lfsr[691], lfsr[692], lfsr[693], lfsr[694], lfsr[695], lfsr[696], lfsr[697], lfsr[698], lfsr[699], lfsr[700], lfsr[701], lfsr[702], lfsr[703], lfsr[704], lfsr[705], lfsr[706], lfsr[707], lfsr[708], lfsr[709], lfsr[710], lfsr[711], lfsr[712], lfsr[713], lfsr[714], lfsr[715], lfsr[716]}; 
//             bits4 <= {lfsr[717], lfsr[718], lfsr[719], lfsr[720], lfsr[721], lfsr[722], lfsr[723], lfsr[724], lfsr[725], lfsr[726], lfsr[727], lfsr[728], lfsr[729], lfsr[730], lfsr[731], lfsr[732], lfsr[733], lfsr[734], lfsr[735], lfsr[736], lfsr[737], lfsr[738], lfsr[739], lfsr[740], lfsr[741], lfsr[742], lfsr[743], lfsr[744], lfsr[745], lfsr[746], lfsr[747], lfsr[748], lfsr[749], lfsr[750], lfsr[751], lfsr[752], lfsr[753], lfsr[754], lfsr[755], lfsr[756], lfsr[757], lfsr[758], lfsr[759], lfsr[760], lfsr[761], lfsr[762], lfsr[763], lfsr[764], lfsr[765], lfsr[766], lfsr[767], lfsr[768], lfsr[769], lfsr[770], lfsr[771], lfsr[772], lfsr[773], lfsr[774], lfsr[775], lfsr[776], lfsr[777], lfsr[778], lfsr[779], lfsr[780], lfsr[781], lfsr[782], lfsr[783], lfsr[784], lfsr[785], lfsr[786], lfsr[787], lfsr[788], lfsr[789], lfsr[790], lfsr[791], lfsr[792], lfsr[793], lfsr[794], lfsr[795], lfsr[796], lfsr[797], lfsr[798], lfsr[799], lfsr[800], lfsr[801], lfsr[802], lfsr[803], lfsr[804], lfsr[805], lfsr[806], lfsr[807], lfsr[808], lfsr[809], lfsr[810], lfsr[811], lfsr[812], lfsr[813], lfsr[814], lfsr[815], lfsr[816], lfsr[817], lfsr[818], lfsr[819], lfsr[820], lfsr[821], lfsr[822], lfsr[823], lfsr[824], lfsr[825], lfsr[826], lfsr[827], lfsr[828], lfsr[829], lfsr[830], lfsr[831], lfsr[832], lfsr[833], lfsr[834], lfsr[835], lfsr[836], lfsr[837], lfsr[838], lfsr[839], lfsr[840], lfsr[841], lfsr[842], lfsr[843], lfsr[844], lfsr[845], lfsr[846], lfsr[847], lfsr[848], lfsr[849], lfsr[850], lfsr[851], lfsr[852], lfsr[853], lfsr[854], lfsr[855], lfsr[856], lfsr[857], lfsr[858], lfsr[859], lfsr[860], lfsr[861], lfsr[862], lfsr[863], lfsr[864], lfsr[865], lfsr[866], lfsr[867], lfsr[868], lfsr[869], lfsr[870], lfsr[871], lfsr[872], lfsr[873], lfsr[874], lfsr[875], lfsr[876], lfsr[877], lfsr[878], lfsr[879], lfsr[880], lfsr[881], lfsr[882], lfsr[883], lfsr[884], lfsr[885], lfsr[886], lfsr[887], lfsr[888], lfsr[889], lfsr[890], lfsr[891], lfsr[892], lfsr[893], lfsr[894], lfsr[895], lfsr[896], lfsr[897], lfsr[898], lfsr[899], lfsr[900], lfsr[901], lfsr[902], lfsr[903], lfsr[904], lfsr[905], lfsr[906], lfsr[907], lfsr[908], lfsr[909], lfsr[910], lfsr[911], lfsr[912], lfsr[913], lfsr[914], lfsr[915], lfsr[916], lfsr[917], lfsr[918], lfsr[919], lfsr[920], lfsr[921], lfsr[922], lfsr[923], lfsr[924], lfsr[925], lfsr[926], lfsr[927], lfsr[928], lfsr[929], lfsr[930], lfsr[931], lfsr[932], lfsr[933], lfsr[934], lfsr[935], lfsr[936], lfsr[937], lfsr[938], lfsr[939], lfsr[940], lfsr[941], lfsr[942], lfsr[943], lfsr[944], lfsr[945], lfsr[946], lfsr[947], lfsr[948], lfsr[949], lfsr[950], lfsr[951], lfsr[952], lfsr[953], lfsr[954], lfsr[955]}; 
//             bits5 <= {lfsr[956], lfsr[957], lfsr[958], lfsr[959], lfsr[960], lfsr[961], lfsr[962], lfsr[963], lfsr[964], lfsr[965], lfsr[966], lfsr[967], lfsr[968], lfsr[969], lfsr[970], lfsr[971], lfsr[972], lfsr[973], lfsr[974], lfsr[975], lfsr[976], lfsr[977], lfsr[978], lfsr[979], lfsr[980], lfsr[981], lfsr[982], lfsr[983], lfsr[984], lfsr[985], lfsr[986], lfsr[987], lfsr[988], lfsr[989], lfsr[990], lfsr[991], lfsr[992], lfsr[993], lfsr[994], lfsr[995], lfsr[996], lfsr[997], lfsr[998], lfsr[999], lfsr[1000], lfsr[1001], lfsr[1002], lfsr[1003], lfsr[1004], lfsr[1005], lfsr[1006], lfsr[1007], lfsr[1008], lfsr[1009], lfsr[1010], lfsr[1011], lfsr[1012], lfsr[1013], lfsr[1014], lfsr[1015], lfsr[1016], lfsr[1017], lfsr[1018], lfsr[1019], lfsr[1020], lfsr[1021], lfsr[1022], lfsr[1023], lfsr[1024], lfsr[1025], lfsr[1026], lfsr[1027], lfsr[1028], lfsr[1029], lfsr[1030], lfsr[1031], lfsr[1032], lfsr[1033], lfsr[1034], lfsr[1035], lfsr[1036], lfsr[1037], lfsr[1038], lfsr[1039], lfsr[1040], lfsr[1041], lfsr[1042], lfsr[1043], lfsr[1044], lfsr[1045], lfsr[1046], lfsr[1047], lfsr[1048], lfsr[1049], lfsr[1050], lfsr[1051], lfsr[1052], lfsr[1053], lfsr[1054], lfsr[1055], lfsr[1056], lfsr[1057], lfsr[1058], lfsr[1059], lfsr[1060], lfsr[1061], lfsr[1062], lfsr[1063], lfsr[1064], lfsr[1065], lfsr[1066], lfsr[1067], lfsr[1068], lfsr[1069], lfsr[1070], lfsr[1071], lfsr[1072], lfsr[1073], lfsr[1074], lfsr[1075], lfsr[1076], lfsr[1077], lfsr[1078], lfsr[1079], lfsr[1080], lfsr[1081], lfsr[1082], lfsr[1083], lfsr[1084], lfsr[1085], lfsr[1086], lfsr[1087], lfsr[1088], lfsr[1089], lfsr[1090], lfsr[1091], lfsr[1092], lfsr[1093], lfsr[1094], lfsr[1095], lfsr[1096], lfsr[1097], lfsr[1098], lfsr[1099], lfsr[1100], lfsr[1101], lfsr[1102], lfsr[1103], lfsr[1104], lfsr[1105], lfsr[1106], lfsr[1107], lfsr[1108], lfsr[1109], lfsr[1110], lfsr[1111], lfsr[1112], lfsr[1113], lfsr[1114], lfsr[1115], lfsr[1116], lfsr[1117], lfsr[1118], lfsr[1119], lfsr[1120], lfsr[1121], lfsr[1122], lfsr[1123], lfsr[1124], lfsr[1125], lfsr[1126], lfsr[1127], lfsr[1128], lfsr[1129], lfsr[1130], lfsr[1131], lfsr[1132], lfsr[1133], lfsr[1134], lfsr[1135], lfsr[1136], lfsr[1137], lfsr[1138], lfsr[1139], lfsr[1140], lfsr[1141], lfsr[1142], lfsr[1143], lfsr[1144], lfsr[1145], lfsr[1146], lfsr[1147], lfsr[1148], lfsr[1149], lfsr[1150], lfsr[1151], lfsr[1152], lfsr[1153], lfsr[1154], lfsr[1155], lfsr[1156], lfsr[1157], lfsr[1158], lfsr[1159], lfsr[1160], lfsr[1161], lfsr[1162], lfsr[1163], lfsr[1164], lfsr[1165], lfsr[1166], lfsr[1167], lfsr[1168], lfsr[1169], lfsr[1170], lfsr[1171], lfsr[1172], lfsr[1173], lfsr[1174], lfsr[1175], lfsr[1176], lfsr[1177], lfsr[1178], lfsr[1179], lfsr[1180], lfsr[1181], lfsr[1182], lfsr[1183], lfsr[1184], lfsr[1185], lfsr[1186], lfsr[1187], lfsr[1188], lfsr[1189], lfsr[1190], lfsr[1191], lfsr[1192], lfsr[1193], lfsr[1194]}; 
//             bits6 <= {lfsr[1195], lfsr[1196], lfsr[1197], lfsr[1198], lfsr[1199], lfsr[1200], lfsr[1201], lfsr[1202], lfsr[1203], lfsr[1204], lfsr[1205], lfsr[1206], lfsr[1207], lfsr[1208], lfsr[1209], lfsr[1210], lfsr[1211], lfsr[1212], lfsr[1213], lfsr[1214], lfsr[1215], lfsr[1216], lfsr[1217], lfsr[1218], lfsr[1219], lfsr[1220], lfsr[1221], lfsr[1222], lfsr[1223], lfsr[1224], lfsr[1225], lfsr[1226], lfsr[1227], lfsr[1228], lfsr[1229], lfsr[1230], lfsr[1231], lfsr[1232], lfsr[1233], lfsr[1234], lfsr[1235], lfsr[1236], lfsr[1237], lfsr[1238], lfsr[1239], lfsr[1240], lfsr[1241], lfsr[1242], lfsr[1243], lfsr[1244], lfsr[1245], lfsr[1246], lfsr[1247], lfsr[1248], lfsr[1249], lfsr[1250], lfsr[1251], lfsr[1252], lfsr[1253], lfsr[1254], lfsr[1255], lfsr[1256], lfsr[1257], lfsr[1258], lfsr[1259], lfsr[1260], lfsr[1261], lfsr[1262], lfsr[1263], lfsr[1264], lfsr[1265], lfsr[1266], lfsr[1267], lfsr[1268], lfsr[1269], lfsr[1270], lfsr[1271], lfsr[1272], lfsr[1273], lfsr[1274], lfsr[1275], lfsr[1276], lfsr[1277], lfsr[1278], lfsr[1279], lfsr[1280], lfsr[1281], lfsr[1282], lfsr[1283], lfsr[1284], lfsr[1285], lfsr[1286], lfsr[1287], lfsr[1288], lfsr[1289], lfsr[1290], lfsr[1291], lfsr[1292], lfsr[1293], lfsr[1294], lfsr[1295], lfsr[1296], lfsr[1297], lfsr[1298], lfsr[1299], lfsr[1300], lfsr[1301], lfsr[1302], lfsr[1303], lfsr[1304], lfsr[1305], lfsr[1306], lfsr[1307], lfsr[1308], lfsr[1309], lfsr[1310], lfsr[1311], lfsr[1312], lfsr[1313], lfsr[1314], lfsr[1315], lfsr[1316], lfsr[1317], lfsr[1318], lfsr[1319], lfsr[1320], lfsr[1321], lfsr[1322], lfsr[1323], lfsr[1324], lfsr[1325], lfsr[1326], lfsr[1327], lfsr[1328], lfsr[1329], lfsr[1330], lfsr[1331], lfsr[1332], lfsr[1333], lfsr[1334], lfsr[1335], lfsr[1336], lfsr[1337], lfsr[1338], lfsr[1339], lfsr[1340], lfsr[1341], lfsr[1342], lfsr[1343], lfsr[1344], lfsr[1345], lfsr[1346], lfsr[1347], lfsr[1348], lfsr[1349], lfsr[1350], lfsr[1351], lfsr[1352], lfsr[1353], lfsr[1354], lfsr[1355], lfsr[1356], lfsr[1357], lfsr[1358], lfsr[1359], lfsr[1360], lfsr[1361], lfsr[1362], lfsr[1363], lfsr[1364], lfsr[1365], lfsr[1366], lfsr[1367], lfsr[1368], lfsr[1369], lfsr[1370], lfsr[1371], lfsr[1372], lfsr[1373], lfsr[1374], lfsr[1375], lfsr[1376], lfsr[1377], lfsr[1378], lfsr[1379], lfsr[1380], lfsr[1381], lfsr[1382], lfsr[1383], lfsr[1384], lfsr[1385], lfsr[1386], lfsr[1387], lfsr[1388], lfsr[1389], lfsr[1390], lfsr[1391], lfsr[1392], lfsr[1393], lfsr[1394], lfsr[1395], lfsr[1396], lfsr[1397], lfsr[1398], lfsr[1399], lfsr[1400], lfsr[1401], lfsr[1402], lfsr[1403], lfsr[1404], lfsr[1405], lfsr[1406], lfsr[1407], lfsr[1408], lfsr[1409], lfsr[1410], lfsr[1411], lfsr[1412], lfsr[1413], lfsr[1414], lfsr[1415], lfsr[1416], lfsr[1417], lfsr[1418], lfsr[1419], lfsr[1420], lfsr[1421], lfsr[1422], lfsr[1423], lfsr[1424], lfsr[1425], lfsr[1426], lfsr[1427], lfsr[1428], lfsr[1429], lfsr[1430], lfsr[1431], lfsr[1432], lfsr[1433]}; 
//             bits7 <= {lfsr[1434], lfsr[1435], lfsr[1436], lfsr[1437], lfsr[1438], lfsr[1439], lfsr[1440], lfsr[1441], lfsr[1442], lfsr[1443], lfsr[1444], lfsr[1445], lfsr[1446], lfsr[1447], lfsr[1448], lfsr[1449], lfsr[1450], lfsr[1451], lfsr[1452], lfsr[1453], lfsr[1454], lfsr[1455], lfsr[1456], lfsr[1457], lfsr[1458], lfsr[1459], lfsr[1460], lfsr[1461], lfsr[1462], lfsr[1463], lfsr[1464], lfsr[1465], lfsr[1466], lfsr[1467], lfsr[1468], lfsr[1469], lfsr[1470], lfsr[1471], lfsr[1472], lfsr[1473], lfsr[1474], lfsr[1475], lfsr[1476], lfsr[1477], lfsr[1478], lfsr[1479], lfsr[1480], lfsr[1481], lfsr[1482], lfsr[1483], lfsr[1484], lfsr[1485], lfsr[1486], lfsr[1487], lfsr[1488], lfsr[1489], lfsr[1490], lfsr[1491], lfsr[1492], lfsr[1493], lfsr[1494], lfsr[1495], lfsr[1496], lfsr[1497], lfsr[1498], lfsr[1499], lfsr[1500], lfsr[1501], lfsr[1502], lfsr[1503], lfsr[1504], lfsr[1505], lfsr[1506], lfsr[1507], lfsr[1508], lfsr[1509], lfsr[1510], lfsr[1511], lfsr[1512], lfsr[1513], lfsr[1514], lfsr[1515], lfsr[1516], lfsr[1517], lfsr[1518], lfsr[1519], lfsr[1520], lfsr[1521], lfsr[1522], lfsr[1523], lfsr[1524], lfsr[1525], lfsr[1526], lfsr[1527], lfsr[1528], lfsr[1529], lfsr[1530], lfsr[1531], lfsr[1532], lfsr[1533], lfsr[1534], lfsr[1535], lfsr[1536], lfsr[1537], lfsr[1538], lfsr[1539], lfsr[1540], lfsr[1541], lfsr[1542], lfsr[1543], lfsr[1544], lfsr[1545], lfsr[1546], lfsr[1547], lfsr[1548], lfsr[1549], lfsr[1550], lfsr[1551], lfsr[1552], lfsr[1553], lfsr[1554], lfsr[1555], lfsr[1556], lfsr[1557], lfsr[1558], lfsr[1559], lfsr[1560], lfsr[1561], lfsr[1562], lfsr[1563], lfsr[1564], lfsr[1565], lfsr[1566], lfsr[1567], lfsr[1568], lfsr[1569], lfsr[1570], lfsr[1571], lfsr[1572], lfsr[1573], lfsr[1574], lfsr[1575], lfsr[1576], lfsr[1577], lfsr[1578], lfsr[1579], lfsr[1580], lfsr[1581], lfsr[1582], lfsr[1583], lfsr[1584], lfsr[1585], lfsr[1586], lfsr[1587], lfsr[1588], lfsr[1589], lfsr[1590], lfsr[1591], lfsr[1592], lfsr[1593], lfsr[1594], lfsr[1595], lfsr[1596], lfsr[1597], lfsr[1598], lfsr[1599], lfsr[1600], lfsr[1601], lfsr[1602], lfsr[1603], lfsr[1604], lfsr[1605], lfsr[1606], lfsr[1607], lfsr[1608], lfsr[1609], lfsr[1610], lfsr[1611], lfsr[1612], lfsr[1613], lfsr[1614], lfsr[1615], lfsr[1616], lfsr[1617], lfsr[1618], lfsr[1619], lfsr[1620], lfsr[1621], lfsr[1622], lfsr[1623], lfsr[1624], lfsr[1625], lfsr[1626], lfsr[1627], lfsr[1628], lfsr[1629], lfsr[1630], lfsr[1631], lfsr[1632], lfsr[1633], lfsr[1634], lfsr[1635], lfsr[1636], lfsr[1637], lfsr[1638], lfsr[1639], lfsr[1640], lfsr[1641], lfsr[1642], lfsr[1643], lfsr[1644], lfsr[1645], lfsr[1646], lfsr[1647], lfsr[1648], lfsr[1649], lfsr[1650], lfsr[1651], lfsr[1652], lfsr[1653], lfsr[1654], lfsr[1655], lfsr[1656], lfsr[1657], lfsr[1658], lfsr[1659], lfsr[1660], lfsr[1661], lfsr[1662], lfsr[1663], lfsr[1664], lfsr[1665], lfsr[1666], lfsr[1667], lfsr[1668], lfsr[1669], lfsr[1670], lfsr[1671], lfsr[1672]}; 
//             bits8 <= {lfsr[1673], lfsr[1674], lfsr[1675], lfsr[1676], lfsr[1677], lfsr[1678], lfsr[1679], lfsr[1680], lfsr[1681], lfsr[1682], lfsr[1683], lfsr[1684], lfsr[1685], lfsr[1686], lfsr[1687], lfsr[1688], lfsr[1689], lfsr[1690], lfsr[1691], lfsr[1692], lfsr[1693], lfsr[1694], lfsr[1695], lfsr[1696], lfsr[1697], lfsr[1698], lfsr[1699], lfsr[1700], lfsr[1701], lfsr[1702], lfsr[1703], lfsr[1704], lfsr[1705], lfsr[1706], lfsr[1707], lfsr[1708], lfsr[1709], lfsr[1710], lfsr[1711], lfsr[1712], lfsr[1713], lfsr[1714], lfsr[1715], lfsr[1716], lfsr[1717], lfsr[1718], lfsr[1719], lfsr[1720], lfsr[1721], lfsr[1722], lfsr[1723], lfsr[1724], lfsr[1725], lfsr[1726], lfsr[1727], lfsr[1728], lfsr[1729], lfsr[1730], lfsr[1731], lfsr[1732], lfsr[1733], lfsr[1734], lfsr[1735], lfsr[1736], lfsr[1737], lfsr[1738], lfsr[1739], lfsr[1740], lfsr[1741], lfsr[1742], lfsr[1743], lfsr[1744], lfsr[1745], lfsr[1746], lfsr[1747], lfsr[1748], lfsr[1749], lfsr[1750], lfsr[1751], lfsr[1752], lfsr[1753], lfsr[1754], lfsr[1755], lfsr[1756], lfsr[1757], lfsr[1758], lfsr[1759], lfsr[1760], lfsr[1761], lfsr[1762], lfsr[1763], lfsr[1764], lfsr[1765], lfsr[1766], lfsr[1767], lfsr[1768], lfsr[1769], lfsr[1770], lfsr[1771], lfsr[1772], lfsr[1773], lfsr[1774], lfsr[1775], lfsr[1776], lfsr[1777], lfsr[1778], lfsr[1779], lfsr[1780], lfsr[1781], lfsr[1782], lfsr[1783], lfsr[1784], lfsr[1785], lfsr[1786], lfsr[1787], lfsr[1788], lfsr[1789], lfsr[1790], lfsr[1791], lfsr[1792], lfsr[1793], lfsr[1794], lfsr[1795], lfsr[1796], lfsr[1797], lfsr[1798], lfsr[1799], lfsr[1800], lfsr[1801], lfsr[1802], lfsr[1803], lfsr[1804], lfsr[1805], lfsr[1806], lfsr[1807], lfsr[1808], lfsr[1809], lfsr[1810], lfsr[1811], lfsr[1812], lfsr[1813], lfsr[1814], lfsr[1815], lfsr[1816], lfsr[1817], lfsr[1818], lfsr[1819], lfsr[1820], lfsr[1821], lfsr[1822], lfsr[1823], lfsr[1824], lfsr[1825], lfsr[1826], lfsr[1827], lfsr[1828], lfsr[1829], lfsr[1830], lfsr[1831], lfsr[1832], lfsr[1833], lfsr[1834], lfsr[1835], lfsr[1836], lfsr[1837], lfsr[1838], lfsr[1839], lfsr[1840], lfsr[1841], lfsr[1842], lfsr[1843], lfsr[1844], lfsr[1845], lfsr[1846], lfsr[1847], lfsr[1848], lfsr[1849], lfsr[1850], lfsr[1851], lfsr[1852], lfsr[1853], lfsr[1854], lfsr[1855], lfsr[1856], lfsr[1857], lfsr[1858], lfsr[1859], lfsr[1860], lfsr[1861], lfsr[1862], lfsr[1863], lfsr[1864], lfsr[1865], lfsr[1866], lfsr[1867], lfsr[1868], lfsr[1869], lfsr[1870], lfsr[1871], lfsr[1872], lfsr[1873], lfsr[1874], lfsr[1875], lfsr[1876], lfsr[1877], lfsr[1878], lfsr[1879], lfsr[1880], lfsr[1881], lfsr[1882], lfsr[1883], lfsr[1884], lfsr[1885], lfsr[1886], lfsr[1887], lfsr[1888], lfsr[1889], lfsr[1890], lfsr[1891], lfsr[1892], lfsr[1893], lfsr[1894], lfsr[1895], lfsr[1896], lfsr[1897], lfsr[1898], lfsr[1899], lfsr[1900], lfsr[1901], lfsr[1902], lfsr[1903], lfsr[1904], lfsr[1905], lfsr[1906], lfsr[1907], lfsr[1908], lfsr[1909], lfsr[1910], lfsr[1911]}; 
//             bits9 <= {lfsr[1912], lfsr[1913], lfsr[1914], lfsr[1915], lfsr[1916], lfsr[1917], lfsr[1918], lfsr[1919], lfsr[1920], lfsr[1921], lfsr[1922], lfsr[1923], lfsr[1924], lfsr[1925], lfsr[1926], lfsr[1927], lfsr[1928], lfsr[1929], lfsr[1930], lfsr[1931], lfsr[1932], lfsr[1933], lfsr[1934], lfsr[1935], lfsr[1936], lfsr[1937], lfsr[1938], lfsr[1939], lfsr[1940], lfsr[1941], lfsr[1942], lfsr[1943], lfsr[1944], lfsr[1945], lfsr[1946], lfsr[1947], lfsr[1948], lfsr[1949], lfsr[1950], lfsr[1951], lfsr[1952], lfsr[1953], lfsr[1954], lfsr[1955], lfsr[1956], lfsr[1957], lfsr[1958], lfsr[1959], lfsr[1960], lfsr[1961], lfsr[1962], lfsr[1963], lfsr[1964], lfsr[1965], lfsr[1966], lfsr[1967], lfsr[1968], lfsr[1969], lfsr[1970], lfsr[1971], lfsr[1972], lfsr[1973], lfsr[1974], lfsr[1975], lfsr[1976], lfsr[1977], lfsr[1978], lfsr[1979], lfsr[1980], lfsr[1981], lfsr[1982], lfsr[1983], lfsr[1984], lfsr[1985], lfsr[1986], lfsr[1987], lfsr[1988], lfsr[1989], lfsr[1990], lfsr[1991], lfsr[1992], lfsr[1993], lfsr[1994], lfsr[1995], lfsr[1996], lfsr[1997], lfsr[1998], lfsr[1999], lfsr[2000], lfsr[2001], lfsr[2002], lfsr[2003], lfsr[2004], lfsr[2005], lfsr[2006], lfsr[2007], lfsr[2008], lfsr[2009], lfsr[2010], lfsr[2011], lfsr[2012], lfsr[2013], lfsr[2014], lfsr[2015], lfsr[2016], lfsr[2017], lfsr[2018], lfsr[2019], lfsr[2020], lfsr[2021], lfsr[2022], lfsr[2023], lfsr[2024], lfsr[2025], lfsr[2026], lfsr[2027], lfsr[2028], lfsr[2029], lfsr[2030], lfsr[2031], lfsr[2032], lfsr[2033], lfsr[2034], lfsr[2035], lfsr[2036], lfsr[2037], lfsr[2038], lfsr[2039], lfsr[2040], lfsr[2041], lfsr[2042], lfsr[2043], lfsr[2044], lfsr[2045], lfsr[2046], lfsr[2047], lfsr[2048], lfsr[2049], lfsr[2050], lfsr[2051], lfsr[2052], lfsr[2053], lfsr[2054], lfsr[2055], lfsr[2056], lfsr[2057], lfsr[2058], lfsr[2059], lfsr[2060], lfsr[2061], lfsr[2062], lfsr[2063], lfsr[2064], lfsr[2065], lfsr[2066], lfsr[2067], lfsr[2068], lfsr[2069], lfsr[2070], lfsr[2071], lfsr[2072], lfsr[2073], lfsr[2074], lfsr[2075], lfsr[2076], lfsr[2077], lfsr[2078], lfsr[2079], lfsr[2080], lfsr[2081], lfsr[2082], lfsr[2083], lfsr[2084], lfsr[2085], lfsr[2086], lfsr[2087], lfsr[2088], lfsr[2089], lfsr[2090], lfsr[2091], lfsr[2092], lfsr[2093], lfsr[2094], lfsr[2095], lfsr[2096], lfsr[2097], lfsr[2098], lfsr[2099], lfsr[2100], lfsr[2101], lfsr[2102], lfsr[2103], lfsr[2104], lfsr[2105], lfsr[2106], lfsr[2107], lfsr[2108], lfsr[2109], lfsr[2110], lfsr[2111], lfsr[2112], lfsr[2113], lfsr[2114], lfsr[2115], lfsr[2116], lfsr[2117], lfsr[2118], lfsr[2119], lfsr[2120], lfsr[2121], lfsr[2122], lfsr[2123], lfsr[2124], lfsr[2125], lfsr[2126], lfsr[2127], lfsr[2128], lfsr[2129], lfsr[2130], lfsr[2131], lfsr[2132], lfsr[2133], lfsr[2134], lfsr[2135], lfsr[2136], lfsr[2137], lfsr[2138], lfsr[2139], lfsr[2140], lfsr[2141], lfsr[2142], lfsr[2143], lfsr[2144], lfsr[2145], lfsr[2146], lfsr[2147], lfsr[2148], lfsr[2149], lfsr[2150]}; 
//             bits10 <= {lfsr[2151], lfsr[2152], lfsr[2153], lfsr[2154], lfsr[2155], lfsr[2156], lfsr[2157], lfsr[2158], lfsr[2159], lfsr[2160], lfsr[2161], lfsr[2162], lfsr[2163], lfsr[2164], lfsr[2165], lfsr[2166], lfsr[2167], lfsr[2168], lfsr[2169], lfsr[2170], lfsr[2171], lfsr[2172], lfsr[2173], lfsr[2174], lfsr[2175], lfsr[2176], lfsr[2177], lfsr[2178], lfsr[2179], lfsr[2180], lfsr[2181], lfsr[2182], lfsr[2183], lfsr[2184], lfsr[2185], lfsr[2186], lfsr[2187], lfsr[2188], lfsr[2189], lfsr[2190], lfsr[2191], lfsr[2192], lfsr[2193], lfsr[2194], lfsr[2195], lfsr[2196], lfsr[2197], lfsr[2198], lfsr[2199], lfsr[2200], lfsr[2201], lfsr[2202], lfsr[2203], lfsr[2204], lfsr[2205], lfsr[2206], lfsr[2207], lfsr[2208], lfsr[2209], lfsr[2210], lfsr[2211], lfsr[2212], lfsr[2213], lfsr[2214], lfsr[2215], lfsr[2216], lfsr[2217], lfsr[2218], lfsr[2219], lfsr[2220], lfsr[2221], lfsr[2222], lfsr[2223], lfsr[2224], lfsr[2225], lfsr[2226], lfsr[2227], lfsr[2228], lfsr[2229], lfsr[2230], lfsr[2231], lfsr[2232], lfsr[2233], lfsr[2234], lfsr[2235], lfsr[2236], lfsr[2237], lfsr[2238], lfsr[2239], lfsr[2240], lfsr[2241], lfsr[2242], lfsr[2243], lfsr[2244], lfsr[2245], lfsr[2246], lfsr[2247], lfsr[2248], lfsr[2249], lfsr[2250], lfsr[2251], lfsr[2252], lfsr[2253], lfsr[2254], lfsr[2255], lfsr[2256], lfsr[2257], lfsr[2258], lfsr[2259], lfsr[2260], lfsr[2261], lfsr[2262], lfsr[2263], lfsr[2264], lfsr[2265], lfsr[2266], lfsr[2267], lfsr[2268], lfsr[2269], lfsr[2270], lfsr[2271], lfsr[2272], lfsr[2273], lfsr[2274], lfsr[2275], lfsr[2276], lfsr[2277], lfsr[2278], lfsr[2279], lfsr[2280], lfsr[2281], lfsr[2282], lfsr[2283], lfsr[2284], lfsr[2285], lfsr[2286], lfsr[2287], lfsr[2288], lfsr[2289], lfsr[2290], lfsr[2291], lfsr[2292], lfsr[2293], lfsr[2294], lfsr[2295], lfsr[2296], lfsr[2297], lfsr[2298], lfsr[2299], lfsr[2300], lfsr[2301], lfsr[2302], lfsr[2303], lfsr[2304], lfsr[2305], lfsr[2306], lfsr[2307], lfsr[2308], lfsr[2309], lfsr[2310], lfsr[2311], lfsr[2312], lfsr[2313], lfsr[2314], lfsr[2315], lfsr[2316], lfsr[2317], lfsr[2318], lfsr[2319], lfsr[2320], lfsr[2321], lfsr[2322], lfsr[2323], lfsr[2324], lfsr[2325], lfsr[2326], lfsr[2327], lfsr[2328], lfsr[2329], lfsr[2330], lfsr[2331], lfsr[2332], lfsr[2333], lfsr[2334], lfsr[2335], lfsr[2336], lfsr[2337], lfsr[2338], lfsr[2339], lfsr[2340], lfsr[2341], lfsr[2342], lfsr[2343], lfsr[2344], lfsr[2345], lfsr[2346], lfsr[2347], lfsr[2348], lfsr[2349], lfsr[2350], lfsr[2351], lfsr[2352], lfsr[2353], lfsr[2354], lfsr[2355], lfsr[2356], lfsr[2357], lfsr[2358], lfsr[2359], lfsr[2360], lfsr[2361], lfsr[2362], lfsr[2363], lfsr[2364], lfsr[2365], lfsr[2366], lfsr[2367], lfsr[2368], lfsr[2369], lfsr[2370], lfsr[2371], lfsr[2372], lfsr[2373], lfsr[2374], lfsr[2375], lfsr[2376], lfsr[2377], lfsr[2378], lfsr[2379], lfsr[2380], lfsr[2381], lfsr[2382], lfsr[2383], lfsr[2384], lfsr[2385], lfsr[2386], lfsr[2387], lfsr[2388], lfsr[2389]}; 
//             bits11 <= {lfsr[2390], lfsr[2391], lfsr[2392], lfsr[2393], lfsr[2394], lfsr[2395], lfsr[2396], lfsr[2397], lfsr[2398], lfsr[2399], lfsr[2400], lfsr[2401], lfsr[2402], lfsr[2403], lfsr[2404], lfsr[2405], lfsr[2406], lfsr[2407], lfsr[2408], lfsr[2409], lfsr[2410], lfsr[2411], lfsr[2412], lfsr[2413], lfsr[2414], lfsr[2415], lfsr[2416], lfsr[2417], lfsr[2418], lfsr[2419], lfsr[2420], lfsr[2421], lfsr[2422], lfsr[2423], lfsr[2424], lfsr[2425], lfsr[2426], lfsr[2427], lfsr[2428], lfsr[2429], lfsr[2430], lfsr[2431], lfsr[2432], lfsr[2433], lfsr[2434], lfsr[2435], lfsr[2436], lfsr[2437], lfsr[2438], lfsr[2439], lfsr[2440], lfsr[2441], lfsr[2442], lfsr[2443], lfsr[2444], lfsr[2445], lfsr[2446], lfsr[2447], lfsr[2448], lfsr[2449], lfsr[2450], lfsr[2451], lfsr[2452], lfsr[2453], lfsr[2454], lfsr[2455], lfsr[2456], lfsr[2457], lfsr[2458], lfsr[2459], lfsr[2460], lfsr[2461], lfsr[2462], lfsr[2463], lfsr[2464], lfsr[2465], lfsr[2466], lfsr[2467], lfsr[2468], lfsr[2469], lfsr[2470], lfsr[2471], lfsr[2472], lfsr[2473], lfsr[2474], lfsr[2475], lfsr[2476], lfsr[2477], lfsr[2478], lfsr[2479], lfsr[2480], lfsr[2481], lfsr[2482], lfsr[2483], lfsr[2484], lfsr[2485], lfsr[2486], lfsr[2487], lfsr[2488], lfsr[2489], lfsr[2490], lfsr[2491], lfsr[2492], lfsr[2493], lfsr[2494], lfsr[2495], lfsr[2496], lfsr[2497], lfsr[2498], lfsr[2499], lfsr[2500], lfsr[2501], lfsr[2502], lfsr[2503], lfsr[2504], lfsr[2505], lfsr[2506], lfsr[2507], lfsr[2508], lfsr[2509], lfsr[2510], lfsr[2511], lfsr[2512], lfsr[2513], lfsr[2514], lfsr[2515], lfsr[2516], lfsr[2517], lfsr[2518], lfsr[2519], lfsr[2520], lfsr[2521], lfsr[2522], lfsr[2523], lfsr[2524], lfsr[2525], lfsr[2526], lfsr[2527], lfsr[2528], lfsr[2529], lfsr[2530], lfsr[2531], lfsr[2532], lfsr[2533], lfsr[2534], lfsr[2535], lfsr[2536], lfsr[2537], lfsr[2538], lfsr[2539], lfsr[2540], lfsr[2541], lfsr[2542], lfsr[2543], lfsr[2544], lfsr[2545], lfsr[2546], lfsr[2547], lfsr[2548], lfsr[2549], lfsr[2550], lfsr[2551], lfsr[2552], lfsr[2553], lfsr[2554], lfsr[2555], lfsr[2556], lfsr[2557], lfsr[2558], lfsr[2559], lfsr[2560], lfsr[2561], lfsr[2562], lfsr[2563], lfsr[2564], lfsr[2565], lfsr[2566], lfsr[2567], lfsr[2568], lfsr[2569], lfsr[2570], lfsr[2571], lfsr[2572], lfsr[2573], lfsr[2574], lfsr[2575], lfsr[2576], lfsr[2577], lfsr[2578], lfsr[2579], lfsr[2580], lfsr[2581], lfsr[2582], lfsr[2583], lfsr[2584], lfsr[2585], lfsr[2586], lfsr[2587], lfsr[2588], lfsr[2589], lfsr[2590], lfsr[2591], lfsr[2592], lfsr[2593], lfsr[2594], lfsr[2595], lfsr[2596], lfsr[2597], lfsr[2598], lfsr[2599], lfsr[2600], lfsr[2601], lfsr[2602], lfsr[2603], lfsr[2604], lfsr[2605], lfsr[2606], lfsr[2607], lfsr[2608], lfsr[2609], lfsr[2610], lfsr[2611], lfsr[2612], lfsr[2613], lfsr[2614], lfsr[2615], lfsr[2616], lfsr[2617], lfsr[2618], lfsr[2619], lfsr[2620], lfsr[2621], lfsr[2622], lfsr[2623], lfsr[2624], lfsr[2625], lfsr[2626], lfsr[2627], lfsr[2628]}; 
//             bits12 <= {lfsr[2629], lfsr[2630], lfsr[2631], lfsr[2632], lfsr[2633], lfsr[2634], lfsr[2635], lfsr[2636], lfsr[2637], lfsr[2638], lfsr[2639], lfsr[2640], lfsr[2641], lfsr[2642], lfsr[2643], lfsr[2644], lfsr[2645], lfsr[2646], lfsr[2647], lfsr[2648], lfsr[2649], lfsr[2650], lfsr[2651], lfsr[2652], lfsr[2653], lfsr[2654], lfsr[2655], lfsr[2656], lfsr[2657], lfsr[2658], lfsr[2659], lfsr[2660], lfsr[2661], lfsr[2662], lfsr[2663], lfsr[2664], lfsr[2665], lfsr[2666], lfsr[2667], lfsr[2668], lfsr[2669], lfsr[2670], lfsr[2671], lfsr[2672], lfsr[2673], lfsr[2674], lfsr[2675], lfsr[2676], lfsr[2677], lfsr[2678], lfsr[2679], lfsr[2680], lfsr[2681], lfsr[2682], lfsr[2683], lfsr[2684], lfsr[2685], lfsr[2686], lfsr[2687], lfsr[2688], lfsr[2689], lfsr[2690], lfsr[2691], lfsr[2692], lfsr[2693], lfsr[2694], lfsr[2695], lfsr[2696], lfsr[2697], lfsr[2698], lfsr[2699], lfsr[2700], lfsr[2701], lfsr[2702], lfsr[2703], lfsr[2704], lfsr[2705], lfsr[2706], lfsr[2707], lfsr[2708], lfsr[2709], lfsr[2710], lfsr[2711], lfsr[2712], lfsr[2713], lfsr[2714], lfsr[2715], lfsr[2716], lfsr[2717], lfsr[2718], lfsr[2719], lfsr[2720], lfsr[2721], lfsr[2722], lfsr[2723], lfsr[2724], lfsr[2725], lfsr[2726], lfsr[2727], lfsr[2728], lfsr[2729], lfsr[2730], lfsr[2731], lfsr[2732], lfsr[2733], lfsr[2734], lfsr[2735], lfsr[2736], lfsr[2737], lfsr[2738], lfsr[2739], lfsr[2740], lfsr[2741], lfsr[2742], lfsr[2743], lfsr[2744], lfsr[2745], lfsr[2746], lfsr[2747], lfsr[2748], lfsr[2749], lfsr[2750], lfsr[2751], lfsr[2752], lfsr[2753], lfsr[2754], lfsr[2755], lfsr[2756], lfsr[2757], lfsr[2758], lfsr[2759], lfsr[2760], lfsr[2761], lfsr[2762], lfsr[2763], lfsr[2764], lfsr[2765], lfsr[2766], lfsr[2767], lfsr[2768], lfsr[2769], lfsr[2770], lfsr[2771], lfsr[2772], lfsr[2773], lfsr[2774], lfsr[2775], lfsr[2776], lfsr[2777], lfsr[2778], lfsr[2779], lfsr[2780], lfsr[2781], lfsr[2782], lfsr[2783], lfsr[2784], lfsr[2785], lfsr[2786], lfsr[2787], lfsr[2788], lfsr[2789], lfsr[2790], lfsr[2791], lfsr[2792], lfsr[2793], lfsr[2794], lfsr[2795], lfsr[2796], lfsr[2797], lfsr[2798], lfsr[2799], lfsr[2800], lfsr[2801], lfsr[2802], lfsr[2803], lfsr[2804], lfsr[2805], lfsr[2806], lfsr[2807], lfsr[2808], lfsr[2809], lfsr[2810], lfsr[2811], lfsr[2812], lfsr[2813], lfsr[2814], lfsr[2815], lfsr[2816], lfsr[2817], lfsr[2818], lfsr[2819], lfsr[2820], lfsr[2821], lfsr[2822], lfsr[2823], lfsr[2824], lfsr[2825], lfsr[2826], lfsr[2827], lfsr[2828], lfsr[2829], lfsr[2830], lfsr[2831], lfsr[2832], lfsr[2833], lfsr[2834], lfsr[2835], lfsr[2836], lfsr[2837], lfsr[2838], lfsr[2839], lfsr[2840], lfsr[2841], lfsr[2842], lfsr[2843], lfsr[2844], lfsr[2845], lfsr[2846], lfsr[2847], lfsr[2848], lfsr[2849], lfsr[2850], lfsr[2851], lfsr[2852], lfsr[2853], lfsr[2854], lfsr[2855], lfsr[2856], lfsr[2857], lfsr[2858], lfsr[2859], lfsr[2860], lfsr[2861], lfsr[2862], lfsr[2863], lfsr[2864], lfsr[2865], lfsr[2866], lfsr[2867]}; 
//             bits13 <= {lfsr[2868], lfsr[2869], lfsr[2870], lfsr[2871], lfsr[2872], lfsr[2873], lfsr[2874], lfsr[2875], lfsr[2876], lfsr[2877], lfsr[2878], lfsr[2879], lfsr[2880], lfsr[2881], lfsr[2882], lfsr[2883], lfsr[2884], lfsr[2885], lfsr[2886], lfsr[2887], lfsr[2888], lfsr[2889], lfsr[2890], lfsr[2891], lfsr[2892], lfsr[2893], lfsr[2894], lfsr[2895], lfsr[2896], lfsr[2897], lfsr[2898], lfsr[2899], lfsr[2900], lfsr[2901], lfsr[2902], lfsr[2903], lfsr[2904], lfsr[2905], lfsr[2906], lfsr[2907], lfsr[2908], lfsr[2909], lfsr[2910], lfsr[2911], lfsr[2912], lfsr[2913], lfsr[2914], lfsr[2915], lfsr[2916], lfsr[2917], lfsr[2918], lfsr[2919], lfsr[2920], lfsr[2921], lfsr[2922], lfsr[2923], lfsr[2924], lfsr[2925], lfsr[2926], lfsr[2927], lfsr[2928], lfsr[2929], lfsr[2930], lfsr[2931], lfsr[2932], lfsr[2933], lfsr[2934], lfsr[2935], lfsr[2936], lfsr[2937], lfsr[2938], lfsr[2939], lfsr[2940], lfsr[2941], lfsr[2942], lfsr[2943], lfsr[2944], lfsr[2945], lfsr[2946], lfsr[2947], lfsr[2948], lfsr[2949], lfsr[2950], lfsr[2951], lfsr[2952], lfsr[2953], lfsr[2954], lfsr[2955], lfsr[2956], lfsr[2957], lfsr[2958], lfsr[2959], lfsr[2960], lfsr[2961], lfsr[2962], lfsr[2963], lfsr[2964], lfsr[2965], lfsr[2966], lfsr[2967], lfsr[2968], lfsr[2969], lfsr[2970], lfsr[2971], lfsr[2972], lfsr[2973], lfsr[2974], lfsr[2975], lfsr[2976], lfsr[2977], lfsr[2978], lfsr[2979], lfsr[2980], lfsr[2981], lfsr[2982], lfsr[2983], lfsr[2984], lfsr[2985], lfsr[2986], lfsr[2987], lfsr[2988], lfsr[2989], lfsr[2990], lfsr[2991], lfsr[2992], lfsr[2993], lfsr[2994], lfsr[2995], lfsr[2996], lfsr[2997], lfsr[2998], lfsr[2999], lfsr[3000], lfsr[3001], lfsr[3002], lfsr[3003], lfsr[3004], lfsr[3005], lfsr[3006], lfsr[3007], lfsr[3008], lfsr[3009], lfsr[3010], lfsr[3011], lfsr[3012], lfsr[3013], lfsr[3014], lfsr[3015], lfsr[3016], lfsr[3017], lfsr[3018], lfsr[3019], lfsr[3020], lfsr[3021], lfsr[3022], lfsr[3023], lfsr[3024], lfsr[3025], lfsr[3026], lfsr[3027], lfsr[3028], lfsr[3029], lfsr[3030], lfsr[3031], lfsr[3032], lfsr[3033], lfsr[3034], lfsr[3035], lfsr[3036], lfsr[3037], lfsr[3038], lfsr[3039], lfsr[3040], lfsr[3041], lfsr[3042], lfsr[3043], lfsr[3044], lfsr[3045], lfsr[3046], lfsr[3047], lfsr[3048], lfsr[3049], lfsr[3050], lfsr[3051], lfsr[3052], lfsr[3053], lfsr[3054], lfsr[3055], lfsr[3056], lfsr[3057], lfsr[3058], lfsr[3059], lfsr[3060], lfsr[3061], lfsr[3062], lfsr[3063], lfsr[3064], lfsr[3065], lfsr[3066], lfsr[3067], lfsr[3068], lfsr[3069], lfsr[3070], lfsr[3071], lfsr[3072], lfsr[3073], lfsr[3074], lfsr[3075], lfsr[3076], lfsr[3077], lfsr[3078], lfsr[3079], lfsr[3080], lfsr[3081], lfsr[3082], lfsr[3083], lfsr[3084], lfsr[3085], lfsr[3086], lfsr[3087], lfsr[3088], lfsr[3089], lfsr[3090], lfsr[3091], lfsr[3092], lfsr[3093], lfsr[3094], lfsr[3095], lfsr[3096], lfsr[3097], lfsr[3098], lfsr[3099], lfsr[3100], lfsr[3101], lfsr[3102], lfsr[3103], lfsr[3104], lfsr[3105], lfsr[3106]}; 
//             bits14 <= {lfsr[3107], lfsr[3108], lfsr[3109], lfsr[3110], lfsr[3111], lfsr[3112], lfsr[3113], lfsr[3114], lfsr[3115], lfsr[3116], lfsr[3117], lfsr[3118], lfsr[3119], lfsr[3120], lfsr[3121], lfsr[3122], lfsr[3123], lfsr[3124], lfsr[3125], lfsr[3126], lfsr[3127], lfsr[3128], lfsr[3129], lfsr[3130], lfsr[3131], lfsr[3132], lfsr[3133], lfsr[3134], lfsr[3135], lfsr[3136], lfsr[3137], lfsr[3138], lfsr[3139], lfsr[3140], lfsr[3141], lfsr[3142], lfsr[3143], lfsr[3144], lfsr[3145], lfsr[3146], lfsr[3147], lfsr[3148], lfsr[3149], lfsr[3150], lfsr[3151], lfsr[3152], lfsr[3153], lfsr[3154], lfsr[3155], lfsr[3156], lfsr[3157], lfsr[3158], lfsr[3159], lfsr[3160], lfsr[3161], lfsr[3162], lfsr[3163], lfsr[3164], lfsr[3165], lfsr[3166], lfsr[3167], lfsr[3168], lfsr[3169], lfsr[3170], lfsr[3171], lfsr[3172], lfsr[3173], lfsr[3174], lfsr[3175], lfsr[3176], lfsr[3177], lfsr[3178], lfsr[3179], lfsr[3180], lfsr[3181], lfsr[3182], lfsr[3183], lfsr[3184], lfsr[3185], lfsr[3186], lfsr[3187], lfsr[3188], lfsr[3189], lfsr[3190], lfsr[3191], lfsr[3192], lfsr[3193], lfsr[3194], lfsr[3195], lfsr[3196], lfsr[3197], lfsr[3198], lfsr[3199], lfsr[3200], lfsr[3201], lfsr[3202], lfsr[3203], lfsr[3204], lfsr[3205], lfsr[3206], lfsr[3207], lfsr[3208], lfsr[3209], lfsr[3210], lfsr[3211], lfsr[3212], lfsr[3213], lfsr[3214], lfsr[3215], lfsr[3216], lfsr[3217], lfsr[3218], lfsr[3219], lfsr[3220], lfsr[3221], lfsr[3222], lfsr[3223], lfsr[3224], lfsr[3225], lfsr[3226], lfsr[3227], lfsr[3228], lfsr[3229], lfsr[3230], lfsr[3231], lfsr[3232], lfsr[3233], lfsr[3234], lfsr[3235], lfsr[3236], lfsr[3237], lfsr[3238], lfsr[3239], lfsr[3240], lfsr[3241], lfsr[3242], lfsr[3243], lfsr[3244], lfsr[3245], lfsr[3246], lfsr[3247], lfsr[3248], lfsr[3249], lfsr[3250], lfsr[3251], lfsr[3252], lfsr[3253], lfsr[3254], lfsr[3255], lfsr[3256], lfsr[3257], lfsr[3258], lfsr[3259], lfsr[3260], lfsr[3261], lfsr[3262], lfsr[3263], lfsr[3264], lfsr[3265], lfsr[3266], lfsr[3267], lfsr[3268], lfsr[3269], lfsr[3270], lfsr[3271], lfsr[3272], lfsr[3273], lfsr[3274], lfsr[3275], lfsr[3276], lfsr[3277], lfsr[3278], lfsr[3279], lfsr[3280], lfsr[3281], lfsr[3282], lfsr[3283], lfsr[3284], lfsr[3285], lfsr[3286], lfsr[3287], lfsr[3288], lfsr[3289], lfsr[3290], lfsr[3291], lfsr[3292], lfsr[3293], lfsr[3294], lfsr[3295], lfsr[3296], lfsr[3297], lfsr[3298], lfsr[3299], lfsr[3300], lfsr[3301], lfsr[3302], lfsr[3303], lfsr[3304], lfsr[3305], lfsr[3306], lfsr[3307], lfsr[3308], lfsr[3309], lfsr[3310], lfsr[3311], lfsr[3312], lfsr[3313], lfsr[3314], lfsr[3315], lfsr[3316], lfsr[3317], lfsr[3318], lfsr[3319], lfsr[3320], lfsr[3321], lfsr[3322], lfsr[3323], lfsr[3324], lfsr[3325], lfsr[3326], lfsr[3327], lfsr[3328], lfsr[3329], lfsr[3330], lfsr[3331], lfsr[3332], lfsr[3333], lfsr[3334], lfsr[3335], lfsr[3336], lfsr[3337], lfsr[3338], lfsr[3339], lfsr[3340], lfsr[3341], lfsr[3342], lfsr[3343], lfsr[3344], lfsr[3345]}; 
//             bits15 <= {lfsr[3346], lfsr[3347], lfsr[3348], lfsr[3349], lfsr[3350], lfsr[3351], lfsr[3352], lfsr[3353], lfsr[3354], lfsr[3355], lfsr[3356], lfsr[3357], lfsr[3358], lfsr[3359], lfsr[3360], lfsr[3361], lfsr[3362], lfsr[3363], lfsr[3364], lfsr[3365], lfsr[3366], lfsr[3367], lfsr[3368], lfsr[3369], lfsr[3370], lfsr[3371], lfsr[3372], lfsr[3373], lfsr[3374], lfsr[3375], lfsr[3376], lfsr[3377], lfsr[3378], lfsr[3379], lfsr[3380], lfsr[3381], lfsr[3382], lfsr[3383], lfsr[3384], lfsr[3385], lfsr[3386], lfsr[3387], lfsr[3388], lfsr[3389], lfsr[3390], lfsr[3391], lfsr[3392], lfsr[3393], lfsr[3394], lfsr[3395], lfsr[3396], lfsr[3397], lfsr[3398], lfsr[3399], lfsr[3400], lfsr[3401], lfsr[3402], lfsr[3403], lfsr[3404], lfsr[3405], lfsr[3406], lfsr[3407], lfsr[3408], lfsr[3409], lfsr[3410], lfsr[3411], lfsr[3412], lfsr[3413], lfsr[3414], lfsr[3415], lfsr[3416], lfsr[3417], lfsr[3418], lfsr[3419], lfsr[3420], lfsr[3421], lfsr[3422], lfsr[3423], lfsr[3424], lfsr[3425], lfsr[3426], lfsr[3427], lfsr[3428], lfsr[3429], lfsr[3430], lfsr[3431], lfsr[3432], lfsr[3433], lfsr[3434], lfsr[3435], lfsr[3436], lfsr[3437], lfsr[3438], lfsr[3439], lfsr[3440], lfsr[3441], lfsr[3442], lfsr[3443], lfsr[3444], lfsr[3445], lfsr[3446], lfsr[3447], lfsr[3448], lfsr[3449], lfsr[3450], lfsr[3451], lfsr[3452], lfsr[3453], lfsr[3454], lfsr[3455], lfsr[3456], lfsr[3457], lfsr[3458], lfsr[3459], lfsr[3460], lfsr[3461], lfsr[3462], lfsr[3463], lfsr[3464], lfsr[3465], lfsr[3466], lfsr[3467], lfsr[3468], lfsr[3469], lfsr[3470], lfsr[3471], lfsr[3472], lfsr[3473], lfsr[3474], lfsr[3475], lfsr[3476], lfsr[3477], lfsr[3478], lfsr[3479], lfsr[3480], lfsr[3481], lfsr[3482], lfsr[3483], lfsr[3484], lfsr[3485], lfsr[3486], lfsr[3487], lfsr[3488], lfsr[3489], lfsr[3490], lfsr[3491], lfsr[3492], lfsr[3493], lfsr[3494], lfsr[3495], lfsr[3496], lfsr[3497], lfsr[3498], lfsr[3499], lfsr[3500], lfsr[3501], lfsr[3502], lfsr[3503], lfsr[3504], lfsr[3505], lfsr[3506], lfsr[3507], lfsr[3508], lfsr[3509], lfsr[3510], lfsr[3511], lfsr[3512], lfsr[3513], lfsr[3514], lfsr[3515], lfsr[3516], lfsr[3517], lfsr[3518], lfsr[3519], lfsr[3520], lfsr[3521], lfsr[3522], lfsr[3523], lfsr[3524], lfsr[3525], lfsr[3526], lfsr[3527], lfsr[3528], lfsr[3529], lfsr[3530], lfsr[3531], lfsr[3532], lfsr[3533], lfsr[3534], lfsr[3535], lfsr[3536], lfsr[3537], lfsr[3538], lfsr[3539], lfsr[3540], lfsr[3541], lfsr[3542], lfsr[3543], lfsr[3544], lfsr[3545], lfsr[3546], lfsr[3547], lfsr[3548], lfsr[3549], lfsr[3550], lfsr[3551], lfsr[3552], lfsr[3553], lfsr[3554], lfsr[3555], lfsr[3556], lfsr[3557], lfsr[3558], lfsr[3559], lfsr[3560], lfsr[3561], lfsr[3562], lfsr[3563], lfsr[3564], lfsr[3565], lfsr[3566], lfsr[3567], lfsr[3568], lfsr[3569], lfsr[3570], lfsr[3571], lfsr[3572], lfsr[3573], lfsr[3574], lfsr[3575], lfsr[3576], lfsr[3577], lfsr[3578], lfsr[3579], lfsr[3580], lfsr[3581], lfsr[3582], lfsr[3583], lfsr[3584]}; 
//             bits16 <= {lfsr[3585], lfsr[3586], lfsr[3587], lfsr[3588], lfsr[3589], lfsr[3590], lfsr[3591], lfsr[3592], lfsr[3593], lfsr[3594], lfsr[3595], lfsr[3596], lfsr[3597], lfsr[3598], lfsr[3599], lfsr[3600], lfsr[3601], lfsr[3602], lfsr[3603], lfsr[3604], lfsr[3605], lfsr[3606], lfsr[3607], lfsr[3608], lfsr[3609], lfsr[3610], lfsr[3611], lfsr[3612], lfsr[3613], lfsr[3614], lfsr[3615], lfsr[3616], lfsr[3617], lfsr[3618], lfsr[3619], lfsr[3620], lfsr[3621], lfsr[3622], lfsr[3623], lfsr[3624], lfsr[3625], lfsr[3626], lfsr[3627], lfsr[3628], lfsr[3629], lfsr[3630], lfsr[3631], lfsr[3632], lfsr[3633], lfsr[3634], lfsr[3635], lfsr[3636], lfsr[3637], lfsr[3638], lfsr[3639], lfsr[3640], lfsr[3641], lfsr[3642], lfsr[3643], lfsr[3644], lfsr[3645], lfsr[3646], lfsr[3647], lfsr[3648], lfsr[3649], lfsr[3650], lfsr[3651], lfsr[3652], lfsr[3653], lfsr[3654], lfsr[3655], lfsr[3656], lfsr[3657], lfsr[3658], lfsr[3659], lfsr[3660], lfsr[3661], lfsr[3662], lfsr[3663], lfsr[3664], lfsr[3665], lfsr[3666], lfsr[3667], lfsr[3668], lfsr[3669], lfsr[3670], lfsr[3671], lfsr[3672], lfsr[3673], lfsr[3674], lfsr[3675], lfsr[3676], lfsr[3677], lfsr[3678], lfsr[3679], lfsr[3680], lfsr[3681], lfsr[3682], lfsr[3683], lfsr[3684], lfsr[3685], lfsr[3686], lfsr[3687], lfsr[3688], lfsr[3689], lfsr[3690], lfsr[3691], lfsr[3692], lfsr[3693], lfsr[3694], lfsr[3695], lfsr[3696], lfsr[3697], lfsr[3698], lfsr[3699], lfsr[3700], lfsr[3701], lfsr[3702], lfsr[3703], lfsr[3704], lfsr[3705], lfsr[3706], lfsr[3707], lfsr[3708], lfsr[3709], lfsr[3710], lfsr[3711], lfsr[3712], lfsr[3713], lfsr[3714], lfsr[3715], lfsr[3716], lfsr[3717], lfsr[3718], lfsr[3719], lfsr[3720], lfsr[3721], lfsr[3722], lfsr[3723], lfsr[3724], lfsr[3725], lfsr[3726], lfsr[3727], lfsr[3728], lfsr[3729], lfsr[3730], lfsr[3731], lfsr[3732], lfsr[3733], lfsr[3734], lfsr[3735], lfsr[3736], lfsr[3737], lfsr[3738], lfsr[3739], lfsr[3740], lfsr[3741], lfsr[3742], lfsr[3743], lfsr[3744], lfsr[3745], lfsr[3746], lfsr[3747], lfsr[3748], lfsr[3749], lfsr[3750], lfsr[3751], lfsr[3752], lfsr[3753], lfsr[3754], lfsr[3755], lfsr[3756], lfsr[3757], lfsr[3758], lfsr[3759], lfsr[3760], lfsr[3761], lfsr[3762], lfsr[3763], lfsr[3764], lfsr[3765], lfsr[3766], lfsr[3767], lfsr[3768], lfsr[3769], lfsr[3770], lfsr[3771], lfsr[3772], lfsr[3773], lfsr[3774], lfsr[3775], lfsr[3776], lfsr[3777], lfsr[3778], lfsr[3779], lfsr[3780], lfsr[3781], lfsr[3782], lfsr[3783], lfsr[3784], lfsr[3785], lfsr[3786], lfsr[3787], lfsr[3788], lfsr[3789], lfsr[3790], lfsr[3791], lfsr[3792], lfsr[3793], lfsr[3794], lfsr[3795], lfsr[3796], lfsr[3797], lfsr[3798], lfsr[3799], lfsr[3800], lfsr[3801], lfsr[3802], lfsr[3803], lfsr[3804], lfsr[3805], lfsr[3806], lfsr[3807], lfsr[3808], lfsr[3809], lfsr[3810], lfsr[3811], lfsr[3812], lfsr[3813], lfsr[3814], lfsr[3815], lfsr[3816], lfsr[3817], lfsr[3818], lfsr[3819], lfsr[3820], lfsr[3821], lfsr[3822], lfsr[3823]}; 

//        end else begin
//             lfsr = seed;
//         end 
//    end