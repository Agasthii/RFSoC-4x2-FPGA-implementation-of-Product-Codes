`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/03/2024 03:03:38 PM
// Design Name: 
// Module Name: bchdecoder_16_7
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bchdecoder_256_239(
    input clk,
    input reset,
    input wire[255:0] r,
    output reg[255:0] dec
    );
    reg [7:0] d; ////////////
    reg d_e;
    
    reg [7:0] S1;
    reg [7:0] S3;

    reg [7:0] sigma0;
    reg [7:0] sigma1;
    reg [7:0] sigma2;


    reg [255:0] r1;
    reg [255:0] r2;
    reg [255:0] r3;
    reg [255:0] r4; ///////////
    reg [255:0] r5; ///////////
    
    reg errs;
    reg errs2;
    reg errs3; ///////////////
    reg errs4; ///////////////
    
    reg [7:0] a0; 
    reg [7:0] a1; 
    reg [7:0] a2; 
    reg [7:0] a3; 
    reg [7:0] a4; 
    reg [7:0] a5; 
    reg [7:0] a6; 
    reg [7:0] a7; 
    reg [7:0] a8; 
    reg [7:0] a9; 
    reg [7:0] a10; 
    reg [7:0] a11; 
    reg [7:0] a12; 
    reg [7:0] a13; 
    reg [7:0] a14; 
    reg [7:0] a15; 
    reg [7:0] a16; 
    reg [7:0] a17; 
    reg [7:0] a18; 
    reg [7:0] a19; 
    reg [7:0] a20; 
    reg [7:0] a21; 
    reg [7:0] a22; 
    reg [7:0] a23; 
    reg [7:0] a24; 
    reg [7:0] a25; 
    reg [7:0] a26; 
    reg [7:0] a27; 
    reg [7:0] a28; 
    reg [7:0] a29; 
    reg [7:0] a30; 
    reg [7:0] a31; 
    reg [7:0] a32; 
    reg [7:0] a33; 
    reg [7:0] a34; 
    reg [7:0] a35; 
    reg [7:0] a36; 
    reg [7:0] a37; 
    reg [7:0] a38; 
    reg [7:0] a39; 
    reg [7:0] a40; 
    reg [7:0] a41; 
    reg [7:0] a42; 
    reg [7:0] a43; 
    reg [7:0] a44; 
    reg [7:0] a45; 
    reg [7:0] a46; 
    reg [7:0] a47; 
    reg [7:0] a48; 
    reg [7:0] a49; 
    reg [7:0] a50; 
    reg [7:0] a51; 
    reg [7:0] a52; 
    reg [7:0] a53; 
    reg [7:0] a54; 
    reg [7:0] a55; 
    reg [7:0] a56; 
    reg [7:0] a57; 
    reg [7:0] a58; 
    reg [7:0] a59; 
    reg [7:0] a60; 
    reg [7:0] a61; 
    reg [7:0] a62; 
    reg [7:0] a63; 
    reg [7:0] a64; 
    reg [7:0] a65; 
    reg [7:0] a66; 
    reg [7:0] a67; 
    reg [7:0] a68; 
    reg [7:0] a69; 
    reg [7:0] a70; 
    reg [7:0] a71; 
    reg [7:0] a72; 
    reg [7:0] a73; 
    reg [7:0] a74; 
    reg [7:0] a75; 
    reg [7:0] a76; 
    reg [7:0] a77; 
    reg [7:0] a78; 
    reg [7:0] a79; 
    reg [7:0] a80; 
    reg [7:0] a81; 
    reg [7:0] a82; 
    reg [7:0] a83; 
    reg [7:0] a84; 
    reg [7:0] a85; 
    reg [7:0] a86; 
    reg [7:0] a87; 
    reg [7:0] a88; 
    reg [7:0] a89; 
    reg [7:0] a90; 
    reg [7:0] a91; 
    reg [7:0] a92; 
    reg [7:0] a93; 
    reg [7:0] a94; 
    reg [7:0] a95; 
    reg [7:0] a96; 
    reg [7:0] a97; 
    reg [7:0] a98; 
    reg [7:0] a99; 
    reg [7:0] a100; 
    reg [7:0] a101; 
    reg [7:0] a102; 
    reg [7:0] a103; 
    reg [7:0] a104; 
    reg [7:0] a105; 
    reg [7:0] a106; 
    reg [7:0] a107; 
    reg [7:0] a108; 
    reg [7:0] a109; 
    reg [7:0] a110; 
    reg [7:0] a111; 
    reg [7:0] a112; 
    reg [7:0] a113; 
    reg [7:0] a114; 
    reg [7:0] a115; 
    reg [7:0] a116; 
    reg [7:0] a117; 
    reg [7:0] a118; 
    reg [7:0] a119; 
    reg [7:0] a120; 
    reg [7:0] a121; 
    reg [7:0] a122; 
    reg [7:0] a123; 
    reg [7:0] a124; 
    reg [7:0] a125; 
    reg [7:0] a126; 
    reg [7:0] a127; 
    reg [7:0] a128; 
    reg [7:0] a129; 
    reg [7:0] a130; 
    reg [7:0] a131; 
    reg [7:0] a132; 
    reg [7:0] a133; 
    reg [7:0] a134; 
    reg [7:0] a135; 
    reg [7:0] a136; 
    reg [7:0] a137; 
    reg [7:0] a138; 
    reg [7:0] a139; 
    reg [7:0] a140; 
    reg [7:0] a141; 
    reg [7:0] a142; 
    reg [7:0] a143; 
    reg [7:0] a144; 
    reg [7:0] a145; 
    reg [7:0] a146; 
    reg [7:0] a147; 
    reg [7:0] a148; 
    reg [7:0] a149; 
    reg [7:0] a150; 
    reg [7:0] a151; 
    reg [7:0] a152; 
    reg [7:0] a153; 
    reg [7:0] a154; 
    reg [7:0] a155; 
    reg [7:0] a156; 
    reg [7:0] a157; 
    reg [7:0] a158; 
    reg [7:0] a159; 
    reg [7:0] a160; 
    reg [7:0] a161; 
    reg [7:0] a162; 
    reg [7:0] a163; 
    reg [7:0] a164; 
    reg [7:0] a165; 
    reg [7:0] a166; 
    reg [7:0] a167; 
    reg [7:0] a168; 
    reg [7:0] a169; 
    reg [7:0] a170; 
    reg [7:0] a171; 
    reg [7:0] a172; 
    reg [7:0] a173; 
    reg [7:0] a174; 
    reg [7:0] a175; 
    reg [7:0] a176; 
    reg [7:0] a177; 
    reg [7:0] a178; 
    reg [7:0] a179; 
    reg [7:0] a180; 
    reg [7:0] a181; 
    reg [7:0] a182; 
    reg [7:0] a183; 
    reg [7:0] a184; 
    reg [7:0] a185; 
    reg [7:0] a186; 
    reg [7:0] a187; 
    reg [7:0] a188; 
    reg [7:0] a189; 
    reg [7:0] a190; 
    reg [7:0] a191; 
    reg [7:0] a192; 
    reg [7:0] a193; 
    reg [7:0] a194; 
    reg [7:0] a195; 
    reg [7:0] a196; 
    reg [7:0] a197; 
    reg [7:0] a198; 
    reg [7:0] a199; 
    reg [7:0] a200; 
    reg [7:0] a201; 
    reg [7:0] a202; 
    reg [7:0] a203; 
    reg [7:0] a204; 
    reg [7:0] a205; 
    reg [7:0] a206; 
    reg [7:0] a207; 
    reg [7:0] a208; 
    reg [7:0] a209; 
    reg [7:0] a210; 
    reg [7:0] a211; 
    reg [7:0] a212; 
    reg [7:0] a213; 
    reg [7:0] a214; 
    reg [7:0] a215; 
    reg [7:0] a216; 
    reg [7:0] a217; 
    reg [7:0] a218; 
    reg [7:0] a219; 
    reg [7:0] a220; 
    reg [7:0] a221; 
    reg [7:0] a222; 
    reg [7:0] a223; 
    reg [7:0] a224; 
    reg [7:0] a225; 
    reg [7:0] a226; 
    reg [7:0] a227; 
    reg [7:0] a228; 
    reg [7:0] a229; 
    reg [7:0] a230; 
    reg [7:0] a231; 
    reg [7:0] a232; 
    reg [7:0] a233; 
    reg [7:0] a234; 
    reg [7:0] a235; 
    reg [7:0] a236; 
    reg [7:0] a237; 
    reg [7:0] a238; 
    reg [7:0] a239; 
    reg [7:0] a240; 
    reg [7:0] a241; 
    reg [7:0] a242; 
    reg [7:0] a243; 
    reg [7:0] a244; 
    reg [7:0] a245; 
    reg [7:0] a246; 
    reg [7:0] a247; 
    reg [7:0] a248; 
    reg [7:0] a249; 
    reg [7:0] a250; 
    reg [7:0] a251; 
    reg [7:0] a252; 
    reg [7:0] a253; 
    reg [7:0] a254;
    
    reg [7:0] a0_1; 
    reg [7:0] a1_1; 
    reg [7:0] a2_1; 
    reg [7:0] a3_1; 
    reg [7:0] a4_1; 
    reg [7:0] a5_1; 
    reg [7:0] a6_1; 
    reg [7:0] a7_1; 
    reg [7:0] a8_1; 
    reg [7:0] a9_1; 
    reg [7:0] a10_1; 
    reg [7:0] a11_1; 
    reg [7:0] a12_1; 
    reg [7:0] a13_1; 
    reg [7:0] a14_1; 
    reg [7:0] a15_1; 
    reg [7:0] a16_1; 
    reg [7:0] a17_1; 
    reg [7:0] a18_1; 
    reg [7:0] a19_1; 
    reg [7:0] a20_1; 
    reg [7:0] a21_1; 
    reg [7:0] a22_1; 
    reg [7:0] a23_1; 
    reg [7:0] a24_1; 
    reg [7:0] a25_1; 
    reg [7:0] a26_1; 
    reg [7:0] a27_1; 
    reg [7:0] a28_1; 
    reg [7:0] a29_1; 
    reg [7:0] a30_1; 
    reg [7:0] a31_1; 
    reg [7:0] a32_1; 
    reg [7:0] a33_1; 
    reg [7:0] a34_1; 
    reg [7:0] a35_1; 
    reg [7:0] a36_1; 
    reg [7:0] a37_1; 
    reg [7:0] a38_1; 
    reg [7:0] a39_1; 
    reg [7:0] a40_1; 
    reg [7:0] a41_1; 
    reg [7:0] a42_1; 
    reg [7:0] a43_1; 
    reg [7:0] a44_1; 
    reg [7:0] a45_1; 
    reg [7:0] a46_1; 
    reg [7:0] a47_1; 
    reg [7:0] a48_1; 
    reg [7:0] a49_1; 
    reg [7:0] a50_1; 
    reg [7:0] a51_1; 
    reg [7:0] a52_1; 
    reg [7:0] a53_1; 
    reg [7:0] a54_1; 
    reg [7:0] a55_1; 
    reg [7:0] a56_1; 
    reg [7:0] a57_1; 
    reg [7:0] a58_1; 
    reg [7:0] a59_1; 
    reg [7:0] a60_1; 
    reg [7:0] a61_1; 
    reg [7:0] a62_1; 
    reg [7:0] a63_1; 
    reg [7:0] a64_1; 
    reg [7:0] a65_1; 
    reg [7:0] a66_1; 
    reg [7:0] a67_1; 
    reg [7:0] a68_1; 
    reg [7:0] a69_1; 
    reg [7:0] a70_1; 
    reg [7:0] a71_1; 
    reg [7:0] a72_1; 
    reg [7:0] a73_1; 
    reg [7:0] a74_1; 
    reg [7:0] a75_1; 
    reg [7:0] a76_1; 
    reg [7:0] a77_1; 
    reg [7:0] a78_1; 
    reg [7:0] a79_1; 
    reg [7:0] a80_1; 
    reg [7:0] a81_1; 
    reg [7:0] a82_1; 
    reg [7:0] a83_1; 
    reg [7:0] a84_1; 
    reg [7:0] a85_1; 
    reg [7:0] a86_1; 
    reg [7:0] a87_1; 
    reg [7:0] a88_1; 
    reg [7:0] a89_1; 
    reg [7:0] a90_1; 
    reg [7:0] a91_1; 
    reg [7:0] a92_1; 
    reg [7:0] a93_1; 
    reg [7:0] a94_1; 
    reg [7:0] a95_1; 
    reg [7:0] a96_1; 
    reg [7:0] a97_1; 
    reg [7:0] a98_1; 
    reg [7:0] a99_1; 
    reg [7:0] a100_1; 
    reg [7:0] a101_1; 
    reg [7:0] a102_1; 
    reg [7:0] a103_1; 
    reg [7:0] a104_1; 
    reg [7:0] a105_1; 
    reg [7:0] a106_1; 
    reg [7:0] a107_1; 
    reg [7:0] a108_1; 
    reg [7:0] a109_1; 
    reg [7:0] a110_1; 
    reg [7:0] a111_1; 
    reg [7:0] a112_1; 
    reg [7:0] a113_1; 
    reg [7:0] a114_1; 
    reg [7:0] a115_1; 
    reg [7:0] a116_1; 
    reg [7:0] a117_1; 
    reg [7:0] a118_1; 
    reg [7:0] a119_1; 
    reg [7:0] a120_1; 
    reg [7:0] a121_1; 
    reg [7:0] a122_1; 
    reg [7:0] a123_1; 
    reg [7:0] a124_1; 
    reg [7:0] a125_1; 
    reg [7:0] a126_1; 
    reg [7:0] a127_1; 
    reg [7:0] a128_1; 
    reg [7:0] a129_1; 
    reg [7:0] a130_1; 
    reg [7:0] a131_1; 
    reg [7:0] a132_1; 
    reg [7:0] a133_1; 
    reg [7:0] a134_1; 
    reg [7:0] a135_1; 
    reg [7:0] a136_1; 
    reg [7:0] a137_1; 
    reg [7:0] a138_1; 
    reg [7:0] a139_1; 
    reg [7:0] a140_1; 
    reg [7:0] a141_1; 
    reg [7:0] a142_1; 
    reg [7:0] a143_1; 
    reg [7:0] a144_1; 
    reg [7:0] a145_1; 
    reg [7:0] a146_1; 
    reg [7:0] a147_1; 
    reg [7:0] a148_1; 
    reg [7:0] a149_1; 
    reg [7:0] a150_1; 
    reg [7:0] a151_1; 
    reg [7:0] a152_1; 
    reg [7:0] a153_1; 
    reg [7:0] a154_1; 
    reg [7:0] a155_1; 
    reg [7:0] a156_1; 
    reg [7:0] a157_1; 
    reg [7:0] a158_1; 
    reg [7:0] a159_1; 
    reg [7:0] a160_1; 
    reg [7:0] a161_1; 
    reg [7:0] a162_1; 
    reg [7:0] a163_1; 
    reg [7:0] a164_1; 
    reg [7:0] a165_1; 
    reg [7:0] a166_1; 
    reg [7:0] a167_1; 
    reg [7:0] a168_1; 
    reg [7:0] a169_1; 
    reg [7:0] a170_1; 
    reg [7:0] a171_1; 
    reg [7:0] a172_1; 
    reg [7:0] a173_1; 
    reg [7:0] a174_1; 
    reg [7:0] a175_1; 
    reg [7:0] a176_1; 
    reg [7:0] a177_1; 
    reg [7:0] a178_1; 
    reg [7:0] a179_1; 
    reg [7:0] a180_1; 
    reg [7:0] a181_1; 
    reg [7:0] a182_1; 
    reg [7:0] a183_1; 
    reg [7:0] a184_1; 
    reg [7:0] a185_1; 
    reg [7:0] a186_1; 
    reg [7:0] a187_1; 
    reg [7:0] a188_1; 
    reg [7:0] a189_1; 
    reg [7:0] a190_1; 
    reg [7:0] a191_1; 
    reg [7:0] a192_1; 
    reg [7:0] a193_1; 
    reg [7:0] a194_1; 
    reg [7:0] a195_1; 
    reg [7:0] a196_1; 
    reg [7:0] a197_1; 
    reg [7:0] a198_1; 
    reg [7:0] a199_1; 
    reg [7:0] a200_1; 
    reg [7:0] a201_1; 
    reg [7:0] a202_1; 
    reg [7:0] a203_1; 
    reg [7:0] a204_1; 
    reg [7:0] a205_1; 
    reg [7:0] a206_1; 
    reg [7:0] a207_1; 
    reg [7:0] a208_1; 
    reg [7:0] a209_1; 
    reg [7:0] a210_1; 
    reg [7:0] a211_1; 
    reg [7:0] a212_1; 
    reg [7:0] a213_1; 
    reg [7:0] a214_1; 
    reg [7:0] a215_1; 
    reg [7:0] a216_1; 
    reg [7:0] a217_1; 
    reg [7:0] a218_1; 
    reg [7:0] a219_1; 
    reg [7:0] a220_1; 
    reg [7:0] a221_1; 
    reg [7:0] a222_1; 
    reg [7:0] a223_1; 
    reg [7:0] a224_1; 
    reg [7:0] a225_1; 
    reg [7:0] a226_1; 
    reg [7:0] a227_1; 
    reg [7:0] a228_1; 
    reg [7:0] a229_1; 
    reg [7:0] a230_1; 
    reg [7:0] a231_1; 
    reg [7:0] a232_1; 
    reg [7:0] a233_1; 
    reg [7:0] a234_1; 
    reg [7:0] a235_1; 
    reg [7:0] a236_1; 
    reg [7:0] a237_1; 
    reg [7:0] a238_1; 
    reg [7:0] a239_1; 
    reg [7:0] a240_1; 
    reg [7:0] a241_1; 
    reg [7:0] a242_1; 
    reg [7:0] a243_1; 
    reg [7:0] a244_1; 
    reg [7:0] a245_1; 
    reg [7:0] a246_1; 
    reg [7:0] a247_1; 
    reg [7:0] a248_1; 
    reg [7:0] a249_1; 
    reg [7:0] a250_1; 
    reg [7:0] a251_1; 
    reg [7:0] a252_1; 
    reg [7:0] a253_1; 
    reg [7:0] a254_1;
    
    reg [7:0] a0_2; 
    reg [7:0] a1_2; 
    reg [7:0] a2_2; 
    reg [7:0] a3_2; 
    reg [7:0] a4_2; 
    reg [7:0] a5_2; 
    reg [7:0] a6_2; 
    reg [7:0] a7_2; 
    reg [7:0] a8_2; 
    reg [7:0] a9_2; 
    reg [7:0] a10_2; 
    reg [7:0] a11_2; 
    reg [7:0] a12_2; 
    reg [7:0] a13_2; 
    reg [7:0] a14_2; 
    reg [7:0] a15_2; 
    reg [7:0] a16_2; 
    reg [7:0] a17_2; 
    reg [7:0] a18_2; 
    reg [7:0] a19_2; 
    reg [7:0] a20_2; 
    reg [7:0] a21_2; 
    reg [7:0] a22_2; 
    reg [7:0] a23_2; 
    reg [7:0] a24_2; 
    reg [7:0] a25_2; 
    reg [7:0] a26_2; 
    reg [7:0] a27_2; 
    reg [7:0] a28_2; 
    reg [7:0] a29_2; 
    reg [7:0] a30_2; 
    reg [7:0] a31_2; 
    reg [7:0] a32_2; 
    reg [7:0] a33_2; 
    reg [7:0] a34_2; 
    reg [7:0] a35_2; 
    reg [7:0] a36_2; 
    reg [7:0] a37_2; 
    reg [7:0] a38_2; 
    reg [7:0] a39_2; 
    reg [7:0] a40_2; 
    reg [7:0] a41_2; 
    reg [7:0] a42_2; 
    reg [7:0] a43_2; 
    reg [7:0] a44_2; 
    reg [7:0] a45_2; 
    reg [7:0] a46_2; 
    reg [7:0] a47_2; 
    reg [7:0] a48_2; 
    reg [7:0] a49_2; 
    reg [7:0] a50_2; 
    reg [7:0] a51_2; 
    reg [7:0] a52_2; 
    reg [7:0] a53_2; 
    reg [7:0] a54_2; 
    reg [7:0] a55_2; 
    reg [7:0] a56_2; 
    reg [7:0] a57_2; 
    reg [7:0] a58_2; 
    reg [7:0] a59_2; 
    reg [7:0] a60_2; 
    reg [7:0] a61_2; 
    reg [7:0] a62_2; 
    reg [7:0] a63_2; 
    reg [7:0] a64_2; 
    reg [7:0] a65_2; 
    reg [7:0] a66_2; 
    reg [7:0] a67_2; 
    reg [7:0] a68_2; 
    reg [7:0] a69_2; 
    reg [7:0] a70_2; 
    reg [7:0] a71_2; 
    reg [7:0] a72_2; 
    reg [7:0] a73_2; 
    reg [7:0] a74_2; 
    reg [7:0] a75_2; 
    reg [7:0] a76_2; 
    reg [7:0] a77_2; 
    reg [7:0] a78_2; 
    reg [7:0] a79_2; 
    reg [7:0] a80_2; 
    reg [7:0] a81_2; 
    reg [7:0] a82_2; 
    reg [7:0] a83_2; 
    reg [7:0] a84_2; 
    reg [7:0] a85_2; 
    reg [7:0] a86_2; 
    reg [7:0] a87_2; 
    reg [7:0] a88_2; 
    reg [7:0] a89_2; 
    reg [7:0] a90_2; 
    reg [7:0] a91_2; 
    reg [7:0] a92_2; 
    reg [7:0] a93_2; 
    reg [7:0] a94_2; 
    reg [7:0] a95_2; 
    reg [7:0] a96_2; 
    reg [7:0] a97_2; 
    reg [7:0] a98_2; 
    reg [7:0] a99_2; 
    reg [7:0] a100_2; 
    reg [7:0] a101_2; 
    reg [7:0] a102_2; 
    reg [7:0] a103_2; 
    reg [7:0] a104_2; 
    reg [7:0] a105_2; 
    reg [7:0] a106_2; 
    reg [7:0] a107_2; 
    reg [7:0] a108_2; 
    reg [7:0] a109_2; 
    reg [7:0] a110_2; 
    reg [7:0] a111_2; 
    reg [7:0] a112_2; 
    reg [7:0] a113_2; 
    reg [7:0] a114_2; 
    reg [7:0] a115_2; 
    reg [7:0] a116_2; 
    reg [7:0] a117_2; 
    reg [7:0] a118_2; 
    reg [7:0] a119_2; 
    reg [7:0] a120_2; 
    reg [7:0] a121_2; 
    reg [7:0] a122_2; 
    reg [7:0] a123_2; 
    reg [7:0] a124_2; 
    reg [7:0] a125_2; 
    reg [7:0] a126_2; 
    reg [7:0] a127_2; 
    reg [7:0] a128_2; 
    reg [7:0] a129_2; 
    reg [7:0] a130_2; 
    reg [7:0] a131_2; 
    reg [7:0] a132_2; 
    reg [7:0] a133_2; 
    reg [7:0] a134_2; 
    reg [7:0] a135_2; 
    reg [7:0] a136_2; 
    reg [7:0] a137_2; 
    reg [7:0] a138_2; 
    reg [7:0] a139_2; 
    reg [7:0] a140_2; 
    reg [7:0] a141_2; 
    reg [7:0] a142_2; 
    reg [7:0] a143_2; 
    reg [7:0] a144_2; 
    reg [7:0] a145_2; 
    reg [7:0] a146_2; 
    reg [7:0] a147_2; 
    reg [7:0] a148_2; 
    reg [7:0] a149_2; 
    reg [7:0] a150_2; 
    reg [7:0] a151_2; 
    reg [7:0] a152_2; 
    reg [7:0] a153_2; 
    reg [7:0] a154_2; 
    reg [7:0] a155_2; 
    reg [7:0] a156_2; 
    reg [7:0] a157_2; 
    reg [7:0] a158_2; 
    reg [7:0] a159_2; 
    reg [7:0] a160_2; 
    reg [7:0] a161_2; 
    reg [7:0] a162_2; 
    reg [7:0] a163_2; 
    reg [7:0] a164_2; 
    reg [7:0] a165_2; 
    reg [7:0] a166_2; 
    reg [7:0] a167_2; 
    reg [7:0] a168_2; 
    reg [7:0] a169_2; 
    reg [7:0] a170_2; 
    reg [7:0] a171_2; 
    reg [7:0] a172_2; 
    reg [7:0] a173_2; 
    reg [7:0] a174_2; 
    reg [7:0] a175_2; 
    reg [7:0] a176_2; 
    reg [7:0] a177_2; 
    reg [7:0] a178_2; 
    reg [7:0] a179_2; 
    reg [7:0] a180_2; 
    reg [7:0] a181_2; 
    reg [7:0] a182_2; 
    reg [7:0] a183_2; 
    reg [7:0] a184_2; 
    reg [7:0] a185_2; 
    reg [7:0] a186_2; 
    reg [7:0] a187_2; 
    reg [7:0] a188_2; 
    reg [7:0] a189_2; 
    reg [7:0] a190_2; 
    reg [7:0] a191_2; 
    reg [7:0] a192_2; 
    reg [7:0] a193_2; 
    reg [7:0] a194_2; 
    reg [7:0] a195_2; 
    reg [7:0] a196_2; 
    reg [7:0] a197_2; 
    reg [7:0] a198_2; 
    reg [7:0] a199_2; 
    reg [7:0] a200_2; 
    reg [7:0] a201_2; 
    reg [7:0] a202_2; 
    reg [7:0] a203_2; 
    reg [7:0] a204_2; 
    reg [7:0] a205_2; 
    reg [7:0] a206_2; 
    reg [7:0] a207_2; 
    reg [7:0] a208_2; 
    reg [7:0] a209_2; 
    reg [7:0] a210_2; 
    reg [7:0] a211_2; 
    reg [7:0] a212_2; 
    reg [7:0] a213_2; 
    reg [7:0] a214_2; 
    reg [7:0] a215_2; 
    reg [7:0] a216_2; 
    reg [7:0] a217_2; 
    reg [7:0] a218_2; 
    reg [7:0] a219_2; 
    reg [7:0] a220_2; 
    reg [7:0] a221_2; 
    reg [7:0] a222_2; 
    reg [7:0] a223_2; 
    reg [7:0] a224_2; 
    reg [7:0] a225_2; 
    reg [7:0] a226_2; 
    reg [7:0] a227_2; 
    reg [7:0] a228_2; 
    reg [7:0] a229_2; 
    reg [7:0] a230_2; 
    reg [7:0] a231_2; 
    reg [7:0] a232_2; 
    reg [7:0] a233_2; 
    reg [7:0] a234_2; 
    reg [7:0] a235_2; 
    reg [7:0] a236_2; 
    reg [7:0] a237_2; 
    reg [7:0] a238_2; 
    reg [7:0] a239_2; 
    reg [7:0] a240_2; 
    reg [7:0] a241_2; 
    reg [7:0] a242_2; 
    reg [7:0] a243_2; 
    reg [7:0] a244_2; 
    reg [7:0] a245_2; 
    reg [7:0] a246_2; 
    reg [7:0] a247_2; 
    reg [7:0] a248_2; 
    reg [7:0] a249_2; 
    reg [7:0] a250_2; 
    reg [7:0] a251_2; 
    reg [7:0] a252_2; 
    reg [7:0] a253_2; 
    reg [7:0] a254_2; 

    
    //////////////////
    reg [254:0] err_vec;
    reg [7:0] temp;
    integer x;
    
    always @(posedge clk) begin
        if(reset) begin
            //Clock cycle 1: Compute syndromes S1 and S3         
            S1[0] <= r[0] ^ r[8] ^ r[12] ^ r[13] ^ r[14] ^ r[18] ^ r[21] ^ r[23] ^ r[24] ^ r[25] ^ r[32] ^ r[33] ^ r[36] ^ r[39] ^ r[42] ^ r[43] ^ r[45] ^ r[46] ^ r[47] ^ r[50] ^ r[56] ^ r[58] ^ r[60] ^ r[61] ^ r[63] ^ r[64] ^ r[66] ^ r[68] ^ r[69] ^ r[72] ^ r[74] ^ r[75] ^ r[80] ^ r[81] ^ r[82] ^ r[83] ^ r[84] ^ r[86] ^ r[87] ^ r[89] ^ r[90] ^ r[91] ^ r[92] ^ r[94] ^ r[96] ^ r[97] ^ r[98] ^ r[100] ^ r[104] ^ r[109] ^ r[110] ^ r[112] ^ r[113] ^ r[117] ^ r[118] ^ r[119] ^ r[120] ^ r[123] ^ r[124] ^ r[125] ^ r[128] ^ r[129] ^ r[133] ^ r[135] ^ r[136] ^ r[138] ^ r[141] ^ r[145] ^ r[147] ^ r[150] ^ r[152] ^ r[154] ^ r[157] ^ r[158] ^ r[159] ^ r[161] ^ r[162] ^ r[163] ^ r[165] ^ r[166] ^ r[169] ^ r[170] ^ r[171] ^ r[172] ^ r[174] ^ r[175] ^ r[176] ^ r[177] ^ r[178] ^ r[179] ^ r[181] ^ r[184] ^ r[185] ^ r[188] ^ r[189] ^ r[191] ^ r[193] ^ r[197] ^ r[198] ^ r[204] ^ r[205] ^ r[206] ^ r[208] ^ r[210] ^ r[212] ^ r[214] ^ r[215] ^ r[216] ^ r[217] ^ r[218] ^ r[221] ^ r[223] ^ r[228] ^ r[231] ^ r[232] ^ r[233] ^ r[234] ^ r[235] ^ r[236] ^ r[237] ^ r[238] ^ r[243] ^ r[245] ^ r[246] ^ r[247] ^ r[248] ^ r[252] ^ r[253];
            S1[1] <= r[1] ^ r[9] ^ r[13] ^ r[14] ^ r[15] ^ r[19] ^ r[22] ^ r[24] ^ r[25] ^ r[26] ^ r[33] ^ r[34] ^ r[37] ^ r[40] ^ r[43] ^ r[44] ^ r[46] ^ r[47] ^ r[48] ^ r[51] ^ r[57] ^ r[59] ^ r[61] ^ r[62] ^ r[64] ^ r[65] ^ r[67] ^ r[69] ^ r[70] ^ r[73] ^ r[75] ^ r[76] ^ r[81] ^ r[82] ^ r[83] ^ r[84] ^ r[85] ^ r[87] ^ r[88] ^ r[90] ^ r[91] ^ r[92] ^ r[93] ^ r[95] ^ r[97] ^ r[98] ^ r[99] ^ r[101] ^ r[105] ^ r[110] ^ r[111] ^ r[113] ^ r[114] ^ r[118] ^ r[119] ^ r[120] ^ r[121] ^ r[124] ^ r[125] ^ r[126] ^ r[129] ^ r[130] ^ r[134] ^ r[136] ^ r[137] ^ r[139] ^ r[142] ^ r[146] ^ r[148] ^ r[151] ^ r[153] ^ r[155] ^ r[158] ^ r[159] ^ r[160] ^ r[162] ^ r[163] ^ r[164] ^ r[166] ^ r[167] ^ r[170] ^ r[171] ^ r[172] ^ r[173] ^ r[175] ^ r[176] ^ r[177] ^ r[178] ^ r[179] ^ r[180] ^ r[182] ^ r[185] ^ r[186] ^ r[189] ^ r[190] ^ r[192] ^ r[194] ^ r[198] ^ r[199] ^ r[205] ^ r[206] ^ r[207] ^ r[209] ^ r[211] ^ r[213] ^ r[215] ^ r[216] ^ r[217] ^ r[218] ^ r[219] ^ r[222] ^ r[224] ^ r[229] ^ r[232] ^ r[233] ^ r[234] ^ r[235] ^ r[236] ^ r[237] ^ r[238] ^ r[239] ^ r[244] ^ r[246] ^ r[247] ^ r[248] ^ r[249] ^ r[253] ^ r[254]; 
            S1[2] <= r[2] ^ r[8] ^ r[10] ^ r[12] ^ r[13] ^ r[15] ^ r[16] ^ r[18] ^ r[20] ^ r[21] ^ r[24] ^ r[26] ^ r[27] ^ r[32] ^ r[33] ^ r[34] ^ r[35] ^ r[36] ^ r[38] ^ r[39] ^ r[41] ^ r[42] ^ r[43] ^ r[44] ^ r[46] ^ r[48] ^ r[49] ^ r[50] ^ r[52] ^ r[56] ^ r[61] ^ r[62] ^ r[64] ^ r[65] ^ r[69] ^ r[70] ^ r[71] ^ r[72] ^ r[75] ^ r[76] ^ r[77] ^ r[80] ^ r[81] ^ r[85] ^ r[87] ^ r[88] ^ r[90] ^ r[93] ^ r[97] ^ r[99] ^ r[102] ^ r[104] ^ r[106] ^ r[109] ^ r[110] ^ r[111] ^ r[113] ^ r[114] ^ r[115] ^ r[117] ^ r[118] ^ r[121] ^ r[122] ^ r[123] ^ r[124] ^ r[126] ^ r[127] ^ r[128] ^ r[129] ^ r[130] ^ r[131] ^ r[133] ^ r[136] ^ r[137] ^ r[140] ^ r[141] ^ r[143] ^ r[145] ^ r[149] ^ r[150] ^ r[156] ^ r[157] ^ r[158] ^ r[160] ^ r[162] ^ r[164] ^ r[166] ^ r[167] ^ r[168] ^ r[169] ^ r[170] ^ r[173] ^ r[175] ^ r[180] ^ r[183] ^ r[184] ^ r[185] ^ r[186] ^ r[187] ^ r[188] ^ r[189] ^ r[190] ^ r[195] ^ r[197] ^ r[198] ^ r[199] ^ r[200] ^ r[204] ^ r[205] ^ r[207] ^ r[215] ^ r[219] ^ r[220] ^ r[221] ^ r[225] ^ r[228] ^ r[230] ^ r[231] ^ r[232] ^ r[239] ^ r[240] ^ r[243] ^ r[246] ^ r[249] ^ r[250] ^ r[252] ^ r[253] ^ r[254];
            S1[3] <= r[3] ^ r[8] ^ r[9] ^ r[11] ^ r[12] ^ r[16] ^ r[17] ^ r[18] ^ r[19] ^ r[22] ^ r[23] ^ r[24] ^ r[27] ^ r[28] ^ r[32] ^ r[34] ^ r[35] ^ r[37] ^ r[40] ^ r[44] ^ r[46] ^ r[49] ^ r[51] ^ r[53] ^ r[56] ^ r[57] ^ r[58] ^ r[60] ^ r[61] ^ r[62] ^ r[64] ^ r[65] ^ r[68] ^ r[69] ^ r[70] ^ r[71] ^ r[73] ^ r[74] ^ r[75] ^ r[76] ^ r[77] ^ r[78] ^ r[80] ^ r[83] ^ r[84] ^ r[87] ^ r[88] ^ r[90] ^ r[92] ^ r[96] ^ r[97] ^ r[103] ^ r[104] ^ r[105] ^ r[107] ^ r[109] ^ r[111] ^ r[113] ^ r[114] ^ r[115] ^ r[116] ^ r[117] ^ r[120] ^ r[122] ^ r[127] ^ r[130] ^ r[131] ^ r[132] ^ r[133] ^ r[134] ^ r[135] ^ r[136] ^ r[137] ^ r[142] ^ r[144] ^ r[145] ^ r[146] ^ r[147] ^ r[151] ^ r[152] ^ r[154] ^ r[162] ^ r[166] ^ r[167] ^ r[168] ^ r[172] ^ r[175] ^ r[177] ^ r[178] ^ r[179] ^ r[186] ^ r[187] ^ r[190] ^ r[193] ^ r[196] ^ r[197] ^ r[199] ^ r[200] ^ r[201] ^ r[204] ^ r[210] ^ r[212] ^ r[214] ^ r[215] ^ r[217] ^ r[218] ^ r[220] ^ r[222] ^ r[223] ^ r[226] ^ r[228] ^ r[229] ^ r[234] ^ r[235] ^ r[236] ^ r[237] ^ r[238] ^ r[240] ^ r[241] ^ r[243] ^ r[244] ^ r[245] ^ r[246] ^ r[248] ^ r[250] ^ r[251] ^ r[252] ^ r[254];
            S1[4] <= r[4] ^ r[8] ^ r[9] ^ r[10] ^ r[14] ^ r[17] ^ r[19] ^ r[20] ^ r[21] ^ r[28] ^ r[29] ^ r[32] ^ r[35] ^ r[38] ^ r[39] ^ r[41] ^ r[42] ^ r[43] ^ r[46] ^ r[52] ^ r[54] ^ r[56] ^ r[57] ^ r[59] ^ r[60] ^ r[62] ^ r[64] ^ r[65] ^ r[68] ^ r[70] ^ r[71] ^ r[76] ^ r[77] ^ r[78] ^ r[79] ^ r[80] ^ r[82] ^ r[83] ^ r[85] ^ r[86] ^ r[87] ^ r[88] ^ r[90] ^ r[92] ^ r[93] ^ r[94] ^ r[96] ^ r[100] ^ r[105] ^ r[106] ^ r[108] ^ r[109] ^ r[113] ^ r[114] ^ r[115] ^ r[116] ^ r[119] ^ r[120] ^ r[121] ^ r[124] ^ r[125] ^ r[129] ^ r[131] ^ r[132] ^ r[134] ^ r[137] ^ r[141] ^ r[143] ^ r[146] ^ r[148] ^ r[150] ^ r[153] ^ r[154] ^ r[155] ^ r[157] ^ r[158] ^ r[159] ^ r[161] ^ r[162] ^ r[165] ^ r[166] ^ r[167] ^ r[168] ^ r[170] ^ r[171] ^ r[172] ^ r[173] ^ r[174] ^ r[175] ^ r[177] ^ r[180] ^ r[181] ^ r[184] ^ r[185] ^ r[187] ^ r[189] ^ r[193] ^ r[194] ^ r[200] ^ r[201] ^ r[202] ^ r[204] ^ r[206] ^ r[208] ^ r[210] ^ r[211] ^ r[212] ^ r[213] ^ r[214] ^ r[217] ^ r[219] ^ r[224] ^ r[227] ^ r[228] ^ r[229] ^ r[230] ^ r[231] ^ r[232] ^ r[233] ^ r[234] ^ r[239] ^ r[241] ^ r[242] ^ r[243] ^ r[244] ^ r[248] ^ r[249] ^ r[251]; 
            S1[5] <= r[5] ^ r[9] ^ r[10] ^ r[11] ^ r[15] ^ r[18] ^ r[20] ^ r[21] ^ r[22] ^ r[29] ^ r[30] ^ r[33] ^ r[36] ^ r[39] ^ r[40] ^ r[42] ^ r[43] ^ r[44] ^ r[47] ^ r[53] ^ r[55] ^ r[57] ^ r[58] ^ r[60] ^ r[61] ^ r[63] ^ r[65] ^ r[66] ^ r[69] ^ r[71] ^ r[72] ^ r[77] ^ r[78] ^ r[79] ^ r[80] ^ r[81] ^ r[83] ^ r[84] ^ r[86] ^ r[87] ^ r[88] ^ r[89] ^ r[91] ^ r[93] ^ r[94] ^ r[95] ^ r[97] ^ r[101] ^ r[106] ^ r[107] ^ r[109] ^ r[110] ^ r[114] ^ r[115] ^ r[116] ^ r[117] ^ r[120] ^ r[121] ^ r[122] ^ r[125] ^ r[126] ^ r[130] ^ r[132] ^ r[133] ^ r[135] ^ r[138] ^ r[142] ^ r[144] ^ r[147] ^ r[149] ^ r[151] ^ r[154] ^ r[155] ^ r[156] ^ r[158] ^ r[159] ^ r[160] ^ r[162] ^ r[163] ^ r[166] ^ r[167] ^ r[168] ^ r[169] ^ r[171] ^ r[172] ^ r[173] ^ r[174] ^ r[175] ^ r[176] ^ r[178] ^ r[181] ^ r[182] ^ r[185] ^ r[186] ^ r[188] ^ r[190] ^ r[194] ^ r[195] ^ r[201] ^ r[202] ^ r[203] ^ r[205] ^ r[207] ^ r[209] ^ r[211] ^ r[212] ^ r[213] ^ r[214] ^ r[215] ^ r[218] ^ r[220] ^ r[225] ^ r[228] ^ r[229] ^ r[230] ^ r[231] ^ r[232] ^ r[233] ^ r[234] ^ r[235] ^ r[240] ^ r[242] ^ r[243] ^ r[244] ^ r[245] ^ r[249] ^ r[250] ^ r[252]; 
            S1[6] <= r[6] ^ r[10] ^ r[11] ^ r[12] ^ r[16] ^ r[19] ^ r[21] ^ r[22] ^ r[23] ^ r[30] ^ r[31] ^ r[34] ^ r[37] ^ r[40] ^ r[41] ^ r[43] ^ r[44] ^ r[45] ^ r[48] ^ r[54] ^ r[56] ^ r[58] ^ r[59] ^ r[61] ^ r[62] ^ r[64] ^ r[66] ^ r[67] ^ r[70] ^ r[72] ^ r[73] ^ r[78] ^ r[79] ^ r[80] ^ r[81] ^ r[82] ^ r[84] ^ r[85] ^ r[87] ^ r[88] ^ r[89] ^ r[90] ^ r[92] ^ r[94] ^ r[95] ^ r[96] ^ r[98] ^ r[102] ^ r[107] ^ r[108] ^ r[110] ^ r[111] ^ r[115] ^ r[116] ^ r[117] ^ r[118] ^ r[121] ^ r[122] ^ r[123] ^ r[126] ^ r[127] ^ r[131] ^ r[133] ^ r[134] ^ r[136] ^ r[139] ^ r[143] ^ r[145] ^ r[148] ^ r[150] ^ r[152] ^ r[155] ^ r[156] ^ r[157] ^ r[159] ^ r[160] ^ r[161] ^ r[163] ^ r[164] ^ r[167] ^ r[168] ^ r[169] ^ r[170] ^ r[172] ^ r[173] ^ r[174] ^ r[175] ^ r[176] ^ r[177] ^ r[179] ^ r[182] ^ r[183] ^ r[186] ^ r[187] ^ r[189] ^ r[191] ^ r[195] ^ r[196] ^ r[202] ^ r[203] ^ r[204] ^ r[206] ^ r[208] ^ r[210] ^ r[212] ^ r[213] ^ r[214] ^ r[215] ^ r[216] ^ r[219] ^ r[221] ^ r[226] ^ r[229] ^ r[230] ^ r[231] ^ r[232] ^ r[233] ^ r[234] ^ r[235] ^ r[236] ^ r[241] ^ r[243] ^ r[244] ^ r[245] ^ r[246] ^ r[250] ^ r[251] ^ r[253]; 
            S1[7] <= r[7] ^ r[11] ^ r[12] ^ r[13] ^ r[17] ^ r[20] ^ r[22] ^ r[23] ^ r[24] ^ r[31] ^ r[32] ^ r[35] ^ r[38] ^ r[41] ^ r[42] ^ r[44] ^ r[45] ^ r[46] ^ r[49] ^ r[55] ^ r[57] ^ r[59] ^ r[60] ^ r[62] ^ r[63] ^ r[65] ^ r[67] ^ r[68] ^ r[71] ^ r[73] ^ r[74] ^ r[79] ^ r[80] ^ r[81] ^ r[82] ^ r[83] ^ r[85] ^ r[86] ^ r[88] ^ r[89] ^ r[90] ^ r[91] ^ r[93] ^ r[95] ^ r[96] ^ r[97] ^ r[99] ^ r[103] ^ r[108] ^ r[109] ^ r[111] ^ r[112] ^ r[116] ^ r[117] ^ r[118] ^ r[119] ^ r[122] ^ r[123] ^ r[124] ^ r[127] ^ r[128] ^ r[132] ^ r[134] ^ r[135] ^ r[137] ^ r[140] ^ r[144] ^ r[146] ^ r[149] ^ r[151] ^ r[153] ^ r[156] ^ r[157] ^ r[158] ^ r[160] ^ r[161] ^ r[162] ^ r[164] ^ r[165] ^ r[168] ^ r[169] ^ r[170] ^ r[171] ^ r[173] ^ r[174] ^ r[175] ^ r[176] ^ r[177] ^ r[178] ^ r[180] ^ r[183] ^ r[184] ^ r[187] ^ r[188] ^ r[190] ^ r[192] ^ r[196] ^ r[197] ^ r[203] ^ r[204] ^ r[205] ^ r[207] ^ r[209] ^ r[211] ^ r[213] ^ r[214] ^ r[215] ^ r[216] ^ r[217] ^ r[220] ^ r[222] ^ r[227] ^ r[230] ^ r[231] ^ r[232] ^ r[233] ^ r[234] ^ r[235] ^ r[236] ^ r[237] ^ r[242] ^ r[244] ^ r[245] ^ r[246] ^ r[247] ^ r[251] ^ r[252] ^ r[254]; 
            
            S3[0] <= r[0] ^ r[4] ^ r[6] ^ r[7] ^ r[8] ^ r[11] ^ r[12] ^ r[13] ^ r[14] ^ r[15] ^ r[20] ^ r[21] ^ r[22] ^ r[23] ^ r[24] ^ r[25] ^ r[27] ^ r[28] ^ r[29] ^ r[30] ^ r[32] ^ r[39] ^ r[40] ^ r[41] ^ r[43] ^ r[45] ^ r[46] ^ r[47] ^ r[49] ^ r[50] ^ r[53] ^ r[54] ^ r[55] ^ r[57] ^ r[58] ^ r[59] ^ r[63] ^ r[66] ^ r[68] ^ r[70] ^ r[72] ^ r[76] ^ r[77] ^ r[78] ^ r[79] ^ r[81] ^ r[82] ^ r[84] ^ r[85] ^ r[89] ^ r[91] ^ r[92] ^ r[93] ^ r[96] ^ r[97] ^ r[98] ^ r[99] ^ r[100] ^ r[105] ^ r[106] ^ r[107] ^ r[108] ^ r[109] ^ r[110] ^ r[112] ^ r[113] ^ r[114] ^ r[115] ^ r[117] ^ r[124] ^ r[125] ^ r[126] ^ r[128] ^ r[130] ^ r[131] ^ r[132] ^ r[134] ^ r[135] ^ r[138] ^ r[139] ^ r[140] ^ r[142] ^ r[143] ^ r[144] ^ r[148] ^ r[151] ^ r[153] ^ r[155] ^ r[157] ^ r[161] ^ r[162] ^ r[163] ^ r[164] ^ r[166] ^ r[167] ^ r[169] ^ r[170] ^ r[174] ^ r[176] ^ r[177] ^ r[178] ^ r[181] ^ r[182] ^ r[183] ^ r[184] ^ r[185] ^ r[190] ^ r[191] ^ r[192] ^ r[193] ^ r[194] ^ r[195] ^ r[197] ^ r[198] ^ r[199] ^ r[200] ^ r[202] ^ r[209] ^ r[210] ^ r[211] ^ r[213] ^ r[215] ^ r[216] ^ r[217] ^ r[219] ^ r[220] ^ r[223] ^ r[224] ^ r[225] ^ r[227] ^ r[228] ^ r[229] ^ r[233] ^ r[236] ^ r[238] ^ r[240] ^ r[242] ^ r[246] ^ r[247] ^ r[248] ^ r[249] ^ r[251] ^ r[252] ^ r[254];
            S3[1] <= r[3] ^ r[5] ^ r[8] ^ r[11] ^ r[16] ^ r[17] ^ r[19] ^ r[23] ^ r[25] ^ r[27] ^ r[28] ^ r[29] ^ r[30] ^ r[31] ^ r[33] ^ r[35] ^ r[37] ^ r[38] ^ r[40] ^ r[42] ^ r[43] ^ r[51] ^ r[53] ^ r[54] ^ r[57] ^ r[59] ^ r[60] ^ r[62] ^ r[63] ^ r[64] ^ r[66] ^ r[69] ^ r[71] ^ r[72] ^ r[73] ^ r[74] ^ r[78] ^ r[79] ^ r[82] ^ r[83] ^ r[88] ^ r[90] ^ r[93] ^ r[96] ^ r[101] ^ r[102] ^ r[104] ^ r[108] ^ r[110] ^ r[112] ^ r[113] ^ r[114] ^ r[115] ^ r[116] ^ r[118] ^ r[120] ^ r[122] ^ r[123] ^ r[125] ^ r[127] ^ r[128] ^ r[136] ^ r[138] ^ r[139] ^ r[142] ^ r[144] ^ r[145] ^ r[147] ^ r[148] ^ r[149] ^ r[151] ^ r[154] ^ r[156] ^ r[157] ^ r[158] ^ r[159] ^ r[163] ^ r[164] ^ r[167] ^ r[168] ^ r[173] ^ r[175] ^ r[178] ^ r[181] ^ r[186] ^ r[187] ^ r[189] ^ r[193] ^ r[195] ^ r[197] ^ r[198] ^ r[199] ^ r[200] ^ r[201] ^ r[203] ^ r[205] ^ r[207] ^ r[208] ^ r[210] ^ r[212] ^ r[213] ^ r[221] ^ r[223] ^ r[224] ^ r[227] ^ r[229] ^ r[230] ^ r[232] ^ r[233] ^ r[234] ^ r[236] ^ r[239] ^ r[241] ^ r[242] ^ r[243] ^ r[244] ^ r[248] ^ r[249] ^ r[252] ^ r[253];
            S3[2] <= r[4] ^ r[5] ^ r[6] ^ r[7] ^ r[8] ^ r[9] ^ r[11] ^ r[12] ^ r[13] ^ r[14] ^ r[16] ^ r[23] ^ r[24] ^ r[25] ^ r[27] ^ r[29] ^ r[30] ^ r[31] ^ r[33] ^ r[34] ^ r[37] ^ r[38] ^ r[39] ^ r[41] ^ r[42] ^ r[43] ^ r[47] ^ r[50] ^ r[52] ^ r[54] ^ r[56] ^ r[60] ^ r[61] ^ r[62] ^ r[63] ^ r[65] ^ r[66] ^ r[68] ^ r[69] ^ r[73] ^ r[75] ^ r[76] ^ r[77] ^ r[80] ^ r[81] ^ r[82] ^ r[83] ^ r[84] ^ r[89] ^ r[90] ^ r[91] ^ r[92] ^ r[93] ^ r[94] ^ r[96] ^ r[97] ^ r[98] ^ r[99] ^ r[101] ^ r[108] ^ r[109] ^ r[110] ^ r[112] ^ r[114] ^ r[115] ^ r[116] ^ r[118] ^ r[119] ^ r[122] ^ r[123] ^ r[124] ^ r[126] ^ r[127] ^ r[128] ^ r[132] ^ r[135] ^ r[137] ^ r[139] ^ r[141] ^ r[145] ^ r[146] ^ r[147] ^ r[148] ^ r[150] ^ r[151] ^ r[153] ^ r[154] ^ r[158] ^ r[160] ^ r[161] ^ r[162] ^ r[165] ^ r[166] ^ r[167] ^ r[168] ^ r[169] ^ r[174] ^ r[175] ^ r[176] ^ r[177] ^ r[178] ^ r[179] ^ r[181] ^ r[182] ^ r[183] ^ r[184] ^ r[186] ^ r[193] ^ r[194] ^ r[195] ^ r[197] ^ r[199] ^ r[200] ^ r[201] ^ r[203] ^ r[204] ^ r[207] ^ r[208] ^ r[209] ^ r[211] ^ r[212] ^ r[213] ^ r[217] ^ r[220] ^ r[222] ^ r[224] ^ r[226] ^ r[230] ^ r[231] ^ r[232] ^ r[233] ^ r[235] ^ r[236] ^ r[238] ^ r[239] ^ r[243] ^ r[245] ^ r[246] ^ r[247] ^ r[250] ^ r[251] ^ r[252] ^ r[253] ^ r[254];
            S3[3] <= r[1] ^ r[3] ^ r[4] ^ r[6] ^ r[8] ^ r[9] ^ r[17] ^ r[19] ^ r[20] ^ r[23] ^ r[25] ^ r[26] ^ r[28] ^ r[29] ^ r[30] ^ r[32] ^ r[35] ^ r[37] ^ r[38] ^ r[39] ^ r[40] ^ r[44] ^ r[45] ^ r[48] ^ r[49] ^ r[54] ^ r[56] ^ r[59] ^ r[62] ^ r[67] ^ r[68] ^ r[70] ^ r[74] ^ r[76] ^ r[78] ^ r[79] ^ r[80] ^ r[81] ^ r[82] ^ r[84] ^ r[86] ^ r[88] ^ r[89] ^ r[91] ^ r[93] ^ r[94] ^ r[102] ^ r[104] ^ r[105] ^ r[108] ^ r[110] ^ r[111] ^ r[113] ^ r[114] ^ r[115] ^ r[117] ^ r[120] ^ r[122] ^ r[123] ^ r[124] ^ r[125] ^ r[129] ^ r[130] ^ r[133] ^ r[134] ^ r[139] ^ r[141] ^ r[144] ^ r[147] ^ r[152] ^ r[153] ^ r[155] ^ r[159] ^ r[161] ^ r[163] ^ r[164] ^ r[165] ^ r[166] ^ r[167] ^ r[169] ^ r[171] ^ r[173] ^ r[174] ^ r[176] ^ r[178] ^ r[179] ^ r[187] ^ r[189] ^ r[190] ^ r[193] ^ r[195] ^ r[196] ^ r[198] ^ r[199] ^ r[200] ^ r[202] ^ r[205] ^ r[207] ^ r[208] ^ r[209] ^ r[210] ^ r[214] ^ r[215] ^ r[218] ^ r[219] ^ r[224] ^ r[226] ^ r[229] ^ r[232] ^ r[237] ^ r[238] ^ r[240] ^ r[244] ^ r[246] ^ r[248] ^ r[249] ^ r[250] ^ r[251] ^ r[252] ^ r[254];
            S3[4] <= r[3] ^ r[7] ^ r[13] ^ r[14] ^ r[18] ^ r[19] ^ r[20] ^ r[26] ^ r[29] ^ r[30] ^ r[31] ^ r[32] ^ r[35] ^ r[36] ^ r[38] ^ r[40] ^ r[43] ^ r[44] ^ r[47] ^ r[50] ^ r[51] ^ r[53] ^ r[54] ^ r[55] ^ r[56] ^ r[57] ^ r[58] ^ r[59] ^ r[60] ^ r[63] ^ r[67] ^ r[68] ^ r[70] ^ r[71] ^ r[73] ^ r[76] ^ r[77] ^ r[78] ^ r[81] ^ r[83] ^ r[88] ^ r[92] ^ r[98] ^ r[99] ^ r[103] ^ r[104] ^ r[105] ^ r[111] ^ r[114] ^ r[115] ^ r[116] ^ r[117] ^ r[120] ^ r[121] ^ r[123] ^ r[125] ^ r[128] ^ r[129] ^ r[132] ^ r[135] ^ r[136] ^ r[138] ^ r[139] ^ r[140] ^ r[141] ^ r[142] ^ r[143] ^ r[144] ^ r[145] ^ r[148] ^ r[152] ^ r[153] ^ r[155] ^ r[156] ^ r[158] ^ r[161] ^ r[162] ^ r[163] ^ r[166] ^ r[168] ^ r[173] ^ r[177] ^ r[183] ^ r[184] ^ r[188] ^ r[189] ^ r[190] ^ r[196] ^ r[199] ^ r[200] ^ r[201] ^ r[202] ^ r[205] ^ r[206] ^ r[208] ^ r[210] ^ r[213] ^ r[214] ^ r[217] ^ r[220] ^ r[221] ^ r[223] ^ r[224] ^ r[225] ^ r[226] ^ r[227] ^ r[228] ^ r[229] ^ r[230] ^ r[233] ^ r[237] ^ r[238] ^ r[240] ^ r[241] ^ r[243] ^ r[246] ^ r[247] ^ r[248] ^ r[251] ^ r[253]; 
            S3[5] <= r[3] ^ r[5] ^ r[6] ^ r[7] ^ r[10] ^ r[11] ^ r[12] ^ r[13] ^ r[14] ^ r[19] ^ r[20] ^ r[21] ^ r[22] ^ r[23] ^ r[24] ^ r[26] ^ r[27] ^ r[28] ^ r[29] ^ r[31] ^ r[38] ^ r[39] ^ r[40] ^ r[42] ^ r[44] ^ r[45] ^ r[46] ^ r[48] ^ r[49] ^ r[52] ^ r[53] ^ r[54] ^ r[56] ^ r[57] ^ r[58] ^ r[62] ^ r[65] ^ r[67] ^ r[69] ^ r[71] ^ r[75] ^ r[76] ^ r[77] ^ r[78] ^ r[80] ^ r[81] ^ r[83] ^ r[84] ^ r[88] ^ r[90] ^ r[91] ^ r[92] ^ r[95] ^ r[96] ^ r[97] ^ r[98] ^ r[99] ^ r[104] ^ r[105] ^ r[106] ^ r[107] ^ r[108] ^ r[109] ^ r[111] ^ r[112] ^ r[113] ^ r[114] ^ r[116] ^ r[123] ^ r[124] ^ r[125] ^ r[127] ^ r[129] ^ r[130] ^ r[131] ^ r[133] ^ r[134] ^ r[137] ^ r[138] ^ r[139] ^ r[141] ^ r[142] ^ r[143] ^ r[147] ^ r[150] ^ r[152] ^ r[154] ^ r[156] ^ r[160] ^ r[161] ^ r[162] ^ r[163] ^ r[165] ^ r[166] ^ r[168] ^ r[169] ^ r[173] ^ r[175] ^ r[176] ^ r[177] ^ r[180] ^ r[181] ^ r[182] ^ r[183] ^ r[184] ^ r[189] ^ r[190] ^ r[191] ^ r[192] ^ r[193] ^ r[194] ^ r[196] ^ r[197] ^ r[198] ^ r[199] ^ r[201] ^ r[208] ^ r[209] ^ r[210] ^ r[212] ^ r[214] ^ r[215] ^ r[216] ^ r[218] ^ r[219] ^ r[222] ^ r[223] ^ r[224] ^ r[226] ^ r[227] ^ r[228] ^ r[232] ^ r[235] ^ r[237] ^ r[239] ^ r[241] ^ r[245] ^ r[246] ^ r[247] ^ r[248] ^ r[250] ^ r[251] ^ r[253] ^ r[254];
            S3[6] <= r[2] ^ r[4] ^ r[7] ^ r[10] ^ r[15] ^ r[16] ^ r[18] ^ r[22] ^ r[24] ^ r[26] ^ r[27] ^ r[28] ^ r[29] ^ r[30] ^ r[32] ^ r[34] ^ r[36] ^ r[37] ^ r[39] ^ r[41] ^ r[42] ^ r[50] ^ r[52] ^ r[53] ^ r[56] ^ r[58] ^ r[59] ^ r[61] ^ r[62] ^ r[63] ^ r[65] ^ r[68] ^ r[70] ^ r[71] ^ r[72] ^ r[73] ^ r[77] ^ r[78] ^ r[81] ^ r[82] ^ r[87] ^ r[89] ^ r[92] ^ r[95] ^ r[100] ^ r[101] ^ r[103] ^ r[107] ^ r[109] ^ r[111] ^ r[112] ^ r[113] ^ r[114] ^ r[115] ^ r[117] ^ r[119] ^ r[121] ^ r[122] ^ r[124] ^ r[126] ^ r[127] ^ r[135] ^ r[137] ^ r[138] ^ r[141] ^ r[143] ^ r[144] ^ r[146] ^ r[147] ^ r[148] ^ r[150] ^ r[153] ^ r[155] ^ r[156] ^ r[157] ^ r[158] ^ r[162] ^ r[163] ^ r[166] ^ r[167] ^ r[172] ^ r[174] ^ r[177] ^ r[180] ^ r[185] ^ r[186] ^ r[188] ^ r[192] ^ r[194] ^ r[196] ^ r[197] ^ r[198] ^ r[199] ^ r[200] ^ r[202] ^ r[204] ^ r[206] ^ r[207] ^ r[209] ^ r[211] ^ r[212] ^ r[220] ^ r[222] ^ r[223] ^ r[226] ^ r[228] ^ r[229] ^ r[231] ^ r[232] ^ r[233] ^ r[235] ^ r[238] ^ r[240] ^ r[241] ^ r[242] ^ r[243] ^ r[247] ^ r[248] ^ r[251] ^ r[252];
            S3[7] <= r[4] ^ r[8] ^ r[14] ^ r[15] ^ r[19] ^ r[20] ^ r[21] ^ r[27] ^ r[30] ^ r[31] ^ r[32] ^ r[33] ^ r[36] ^ r[37] ^ r[39] ^ r[41] ^ r[44] ^ r[45] ^ r[48] ^ r[51] ^ r[52] ^ r[54] ^ r[55] ^ r[56] ^ r[57] ^ r[58] ^ r[59] ^ r[60] ^ r[61] ^ r[64] ^ r[68] ^ r[69] ^ r[71] ^ r[72] ^ r[74] ^ r[77] ^ r[78] ^ r[79] ^ r[82] ^ r[84] ^ r[89] ^ r[93] ^ r[99] ^ r[100] ^ r[104] ^ r[105] ^ r[106] ^ r[112] ^ r[115] ^ r[116] ^ r[117] ^ r[118] ^ r[121] ^ r[122] ^ r[124] ^ r[126] ^ r[129] ^ r[130] ^ r[133] ^ r[136] ^ r[137] ^ r[139] ^ r[140] ^ r[141] ^ r[142] ^ r[143] ^ r[144] ^ r[145] ^ r[146] ^ r[149] ^ r[153] ^ r[154] ^ r[156] ^ r[157] ^ r[159] ^ r[162] ^ r[163] ^ r[164] ^ r[167] ^ r[169] ^ r[174] ^ r[178] ^ r[184] ^ r[185] ^ r[189] ^ r[190] ^ r[191] ^ r[197] ^ r[200] ^ r[201] ^ r[202] ^ r[203] ^ r[206] ^ r[207] ^ r[209] ^ r[211] ^ r[214] ^ r[215] ^ r[218] ^ r[221] ^ r[222] ^ r[224] ^ r[225] ^ r[226] ^ r[227] ^ r[228] ^ r[229] ^ r[230] ^ r[231] ^ r[234] ^ r[238] ^ r[239] ^ r[241] ^ r[242] ^ r[244] ^ r[247] ^ r[248] ^ r[249] ^ r[252] ^ r[254];
           
            r1 <= r;
        
            //Clock cycle 2: Compute coefficients of the Peterson Equation    
            sigma0[0] <= S3[0] ^ S1[0] ^ S1[7] ^ S1[4] ^ S1[6] ^ (S1[0] & S1[4]) ^ (S1[0] & S1[6]) ^ (S1[0] & S1[7]) ^ (S1[4] & S1[6]) ^ (S1[2] & S1[4]) ^ (S1[7] & S1[4]) ^ (S1[5] & S1[3]) ^ (S1[3] & S1[7]) ^ (S1[3] & S1[2]) ^ (S1[3] & S1[6]) ^ (S1[5] & S1[2]) ^ (S1[6] & S1[2]);
            sigma0[1] <= S3[1] ^ S1[3] ^ S1[5] ^ (S1[0] & S1[1]) ^ (S1[4] & S1[1]) ^ (S1[6] & S1[1]) ^ (S1[7] & S1[0]) ^ (S1[4] & S1[7]) ^ (S1[4] & S1[6]) ^ (S1[2] & S1[5]) ^ (S1[3] & S1[7]) ^ (S1[5] & S1[3]) ^ (S1[5] & S1[7]) ^ (S1[6] & S1[3]) ^ (S1[6] & S1[7]) ^ (S1[6] & S1[2]);
            sigma0[2] <= S3[2] ^ S1[4] ^ S1[5] ^ S1[6] ^ S1[7] ^ (S1[7] & S1[2]) ^ (S1[0] & S1[1]) ^ (S1[0] & S1[4]) ^ (S1[0] & S1[5]) ^ (S1[0] & S1[6]) ^ (S1[4] & S1[5]) ^ (S1[7] & S1[6]) ^ (S1[5] & S1[3]) ^ (S1[3] & S1[2]) ^ (S1[5] & S1[2]) ^ (S1[6] & S1[4]) ^ (S1[6] & S1[5]) ^ (S1[2] & S1[0]) ^ (S1[1] & S1[7]) ^ (S1[4] & S1[3]) ^ (S1[6] & S1[2]) ^ (S1[7] & S1[3]);
//            sigma0[2] <= S3[2] ^ S1[4] ^ S1[5] ^ S1[6] ^ S1[7] ^ (S1[0] & S1[3]) ^ (S1[7] & S1[2]) ^ (S1[0] & S1[1]) ^ (S1[0] & S1[4]) ^ (S1[0] & S1[5]) ^ (S1[0] & S1[6]) ^ (S1[4] & S1[5]) ^ (S1[2] & S1[4]) ^ (S1[7] & S1[6]) ^ (S1[5] & S1[3]) ^ (S1[3] & S1[2]) ^ (S1[5] & S1[2]) ^ (S1[6] & S1[4]) ^ (S1[3] & S1[6]) ^ (S1[6] & S1[5]);
            sigma0[3] <= S3[3] ^ S1[1] ^ S1[3] ^ S1[4] ^ S1[6] ^ (S1[0] & S1[4]) ^ (S1[0] & S1[6]) ^ (S1[1] & S1[4]) ^ (S1[1] & S1[5]) ^ (S1[2] & S1[3]) ^ (S1[3] & S1[0]) ^ (S1[4] & S1[3]) ^ (S1[3] & S1[7]) ^ (S1[4] & S1[2]) ^ (S1[5] & S1[3]) ^ (S1[6] & S1[1]) ^ (S1[6] & S1[4]) ^ (S1[6] & S1[3]) ^ (S1[7] & S1[1]) ^ (S1[7] & S1[6]) ^ (S1[7] & S1[4]);
            sigma0[4] <= S3[4] ^ S1[3] ^ S1[7] ^ (S1[0] & S1[2]) ^ (S1[0] & S1[5]) ^ (S1[0] & S1[7]) ^ (S1[1] & S1[4]) ^ (S1[2] & S1[1]) ^ (S1[2] & S1[3]) ^ (S1[3] & S1[7]) ^ (S1[4] & S1[3]) ^ (S1[5] & S1[4]) ^ (S1[5] & S1[2]) ^ (S1[6] & S1[1]) ^ (S1[6] & S1[4]) ^ (S1[6] & S1[5]) ^ (S1[7] & S1[1]);
            sigma0[5] <= S3[5] ^ S1[3] ^ S1[5] ^ S1[6] ^ S1[7] ^ (S1[1] & S1[2]) ^ (S1[1] & S1[4]) ^ (S1[1] & S1[5]) ^ (S1[2] & S1[4]) ^ (S1[3] & S1[1]) ^ (S1[3] & S1[6]) ^ (S1[5] & S1[2]) ^ (S1[5] & S1[3]) ^ (S1[6] & S1[2]) ^ (S1[7] & S1[6]) ^ (S1[7] & S1[2]);
            sigma0[6] <= S3[6] ^ S1[2] ^ S1[4] ^ S1[7] ^ (S1[0] & S1[3]) ^ (S1[0] & S1[5]) ^ (S1[1] & S1[5]) ^ (S1[2] & S1[4]) ^ (S1[2] & S1[5]) ^ (S1[4] & S1[1]) ^ (S1[4] & S1[6]) ^ (S1[5] & S1[7]) ^ (S1[5] & S1[3]) ^ (S1[6] & S1[2]) ^ (S1[6] & S1[5]) ^ (S1[6] & S1[3]) ^ (S1[7] & S1[6]);
            sigma0[7] <= S3[7] ^ S1[4] ^ (S1[0] & S1[6]) ^ (S1[1] & S1[3]) ^ (S1[1] & S1[6]) ^ (S1[2] & S1[5]) ^ (S1[3] & S1[2]) ^ (S1[3] & S1[4]) ^ (S1[5] & S1[4]) ^ (S1[5] & S1[6]) ^ (S1[6] & S1[7]) ^ (S1[6] & S1[3]) ^ (S1[7] & S1[0]) ^ (S1[7] & S1[2]) ^ (S1[7] & S1[5]);
            
            
            
            sigma1[0] <= S1[0] ^ S1[4] ^ S1[6] ^ S1[7];
            sigma1[1] <= S1[7];
            sigma1[2] <= S1[1] ^ S1[4] ^ S1[5] ^ S1[6];
            sigma1[3] <= S1[4] ^ S1[6];
            sigma1[4] <= S1[2] ^ S1[4] ^ S1[5] ^ S1[7];
            sigma1[5] <= S1[5];
            sigma1[6] <= S1[3] ^ S1[5] ^ S1[6];
            sigma1[7] <= S1[6];
            
            sigma2 <= S1;
            errs <= !((S1 == 8'b0) & (S3 == 8'b0));
            r2 <= r1;

            
            //Clock cycle 3: Chien Search 
            a0 <= sigma0 ^ sigma1 ^ sigma2; 
            a1 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]); 
            a2 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a3 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a4 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a5 <= sigma0 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a6 <= sigma0 ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a7 <= sigma0 ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a8 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a9 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a10 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a11 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a12 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a13 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]); 
            a14 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a15 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a16 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a17 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a18 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a19 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a20 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a21 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a22 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a23 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a24 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a25 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]); 
            a26 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a27 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a28 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a29 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a30 <= sigma0 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a31 <= sigma0 ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a32 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a33 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a34 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a35 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a36 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a37 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a38 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a39 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a40 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a41 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a42 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a43 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a44 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a45 <= sigma0 ^ sigma1 ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a46 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a47 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a48 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a49 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a50 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a51 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a52 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a53 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a54 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a55 <= sigma0 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a56 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a57 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a58 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a59 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a60 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a61 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a62 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a63 <= sigma0 ^ sigma1 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a64 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a65 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a66 <= sigma0 ^ sigma1 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a67 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a68 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a69 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a70 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a71 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a72 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a73 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a74 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a75 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a76 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a77 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a78 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a79 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a80 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a81 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a82 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a83 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a84 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a85 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a86 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a87 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a88 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a89 <= sigma0 ^ sigma1 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a90 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a91 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a92 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a93 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a94 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a95 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a96 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a97 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a98 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a99 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]); 
            a100 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a101 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a102 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a103 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a104 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a105 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a106 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a107 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a108 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a109 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a110 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a111 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a112 <= sigma0 ^ sigma1 ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a113 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a114 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a115 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a116 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a117 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a118 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a119 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a120 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a121 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a122 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a123 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a124 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a125 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a126 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a127 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a128 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]); 
            a129 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a130 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a131 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a132 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a133 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a134 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a135 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a136 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a137 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a138 <= sigma0 ^ sigma1 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a139 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a140 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]); 
            a141 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a142 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a143 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a144 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a145 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a146 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a147 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a148 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a149 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a150 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a151 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a152 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a153 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a154 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a155 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a156 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a157 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a158 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a159 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a160 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a161 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a162 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a163 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a164 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a165 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a166 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a167 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a168 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a169 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a170 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a171 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a172 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a173 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a174 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a175 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a176 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a177 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a178 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a179 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a180 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a181 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a182 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a183 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a184 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a185 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a186 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a187 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a188 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a189 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a190 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a191 <= sigma0 ^ sigma1 ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a192 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a193 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a194 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a195 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a196 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a197 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a198 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a199 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a200 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a201 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a202 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a203 <= sigma0 ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a204 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a205 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a206 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a207 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a208 <= sigma0 ^ sigma1 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a209 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a210 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a211 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a212 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a213 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a214 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a215 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a216 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a217 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a218 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a219 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a220 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a221 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a222 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a223 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ sigma2 ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a224 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a225 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a226 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a227 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a228 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a229 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a230 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a231 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a232 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a233 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a234 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a235 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a236 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a237 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a238 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a239 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]); 
            a240 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a241 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a242 <= sigma0 ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a243 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a244 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a245 <= sigma0 ^ sigma1 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a246 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a247 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]); 
            a248 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a249 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ sigma2 ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
            a250 <= sigma0 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ sigma2 ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a251 <= sigma0 ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<4) ^ (8'd29 * sigma1[4]) ^ (8'd58 * sigma1[5]) ^ (8'd116 * sigma1[6]) ^ (8'd232 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a252 <= sigma0 ^ sigma1 ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<5) ^ (8'd29 * sigma1[3]) ^ (8'd58 * sigma1[4]) ^ (8'd116 * sigma1[5]) ^ (8'd232 * sigma1[6]) ^ (8'd205 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<5) ^ (8'd29 * sigma2[3]) ^ (8'd58 * sigma2[4]) ^ (8'd116 * sigma2[5]) ^ (8'd232 * sigma2[6]) ^ (8'd205 * sigma2[7]); 
            a253 <= sigma0 ^ sigma1 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<6) ^ (8'd29 * sigma1[2]) ^ (8'd58 * sigma1[3]) ^ (8'd116 * sigma1[4]) ^ (8'd232 * sigma1[5]) ^ (8'd205 * sigma1[6]) ^ (8'd135 * sigma1[7]) ^ (sigma2<<3) ^ (8'd29 * sigma2[5]) ^ (8'd58 * sigma2[6]) ^ (8'd116 * sigma2[7]) ^ (sigma2<<4) ^ (8'd29 * sigma2[4]) ^ (8'd58 * sigma2[5]) ^ (8'd116 * sigma2[6]) ^ (8'd232 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]) ^ (sigma2<<7) ^ (8'd29 * sigma2[1]) ^ (8'd58 * sigma2[2]) ^ (8'd116 * sigma2[3]) ^ (8'd232 * sigma2[4]) ^ (8'd205 * sigma2[5]) ^ (8'd135 * sigma2[6]) ^ (8'd19 * sigma2[7]); 
            a254 <= sigma0 ^ (sigma1<<1) ^ (8'd29 * sigma1[7]) ^ (sigma1<<2) ^ (8'd29 * sigma1[6]) ^ (8'd58 * sigma1[7]) ^ (sigma1<<3) ^ (8'd29 * sigma1[5]) ^ (8'd58 * sigma1[6]) ^ (8'd116 * sigma1[7]) ^ (sigma1<<7) ^ (8'd29 * sigma1[1]) ^ (8'd58 * sigma1[2]) ^ (8'd116 * sigma1[3]) ^ (8'd232 * sigma1[4]) ^ (8'd205 * sigma1[5]) ^ (8'd135 * sigma1[6]) ^ (8'd19 * sigma1[7]) ^ sigma2 ^ (sigma2<<1) ^ (8'd29 * sigma2[7]) ^ (sigma2<<2) ^ (8'd29 * sigma2[6]) ^ (8'd58 * sigma2[7]) ^ (sigma2<<6) ^ (8'd29 * sigma2[2]) ^ (8'd58 * sigma2[3]) ^ (8'd116 * sigma2[4]) ^ (8'd232 * sigma2[5]) ^ (8'd205 * sigma2[6]) ^ (8'd135 * sigma2[7]); 
 
 
            
            
            errs2 <= errs;
            r3 <= r2;
//            d_e <= (|sigma0) ^ (^r2);
//            d <= |sigma0;
            
            //Clock Cycle 4: Error vector
            
            err_vec[0]  <= (a0  == 8'b0) & errs2 ? 1 : 0;
            err_vec[1]  <= (a1  == 8'b0) & errs2 ? 1 : 0;
            err_vec[2]  <= (a2  == 8'b0) & errs2 ? 1 : 0;
            err_vec[3]  <= (a3  == 8'b0) & errs2 ? 1 : 0;
            err_vec[4]  <= (a4  == 8'b0) & errs2 ? 1 : 0;
            err_vec[5]  <= (a5  == 8'b0) & errs2 ? 1 : 0;
            err_vec[6]  <= (a6  == 8'b0) & errs2 ? 1 : 0;
            err_vec[7]  <= (a7  == 8'b0) & errs2 ? 1 : 0;
            err_vec[8]  <= (a8  == 8'b0) & errs2 ? 1 : 0;
            err_vec[9]  <= (a9  == 8'b0) & errs2 ? 1 : 0;
            err_vec[10] <= (a10 == 8'b0) & errs2 ? 1 : 0;
            err_vec[11] <= (a11 == 8'b0) & errs2 ? 1 : 0;
            err_vec[12] <= (a12 == 8'b0) & errs2 ? 1 : 0;
            err_vec[13] <= (a13 == 8'b0) & errs2 ? 1 : 0;
            err_vec[14] <= (a14 == 8'b0) & errs2 ? 1 : 0;
            err_vec[15] <= (a15 == 8'b0) & errs2 ? 1 : 0;
            err_vec[16] <= (a16 == 8'b0) & errs2 ? 1 : 0;
            err_vec[17] <= (a17 == 8'b0) & errs2 ? 1 : 0;
            err_vec[18] <= (a18 == 8'b0) & errs2 ? 1 : 0;
            err_vec[19] <= (a19 == 8'b0) & errs2 ? 1 : 0;
            err_vec[20] <= (a20 == 8'b0) & errs2 ? 1 : 0;
            err_vec[21] <= (a21 == 8'b0) & errs2 ? 1 : 0;
            err_vec[22] <= (a22 == 8'b0) & errs2 ? 1 : 0;
            err_vec[23] <= (a23 == 8'b0) & errs2 ? 1 : 0;
            err_vec[24] <= (a24 == 8'b0) & errs2 ? 1 : 0;
            err_vec[25] <= (a25 == 8'b0) & errs2 ? 1 : 0;
            err_vec[26] <= (a26 == 8'b0) & errs2 ? 1 : 0;
            err_vec[27] <= (a27 == 8'b0) & errs2 ? 1 : 0;
            err_vec[28] <= (a28 == 8'b0) & errs2 ? 1 : 0;
            err_vec[29] <= (a29 == 8'b0) & errs2 ? 1 : 0;
            err_vec[30] <= (a30 == 8'b0) & errs2 ? 1 : 0;
            err_vec[31] <= (a31 == 8'b0) & errs2 ? 1 : 0;
            err_vec[32] <= (a32 == 8'b0) & errs2 ? 1 : 0;
            err_vec[33] <= (a33 == 8'b0) & errs2 ? 1 : 0;
            err_vec[34] <= (a34 == 8'b0) & errs2 ? 1 : 0;
            err_vec[35] <= (a35 == 8'b0) & errs2 ? 1 : 0;
            err_vec[36] <= (a36 == 8'b0) & errs2 ? 1 : 0;
            err_vec[37] <= (a37 == 8'b0) & errs2 ? 1 : 0;
            err_vec[38] <= (a38 == 8'b0) & errs2 ? 1 : 0;
            err_vec[39] <= (a39 == 8'b0) & errs2 ? 1 : 0;
            err_vec[40] <= (a40 == 8'b0) & errs2 ? 1 : 0;
            err_vec[41] <= (a41 == 8'b0) & errs2 ? 1 : 0;
            err_vec[42] <= (a42 == 8'b0) & errs2 ? 1 : 0;
            err_vec[43] <= (a43 == 8'b0) & errs2 ? 1 : 0;
            err_vec[44] <= (a44 == 8'b0) & errs2 ? 1 : 0;
            err_vec[45] <= (a45 == 8'b0) & errs2 ? 1 : 0;
            err_vec[46] <= (a46 == 8'b0) & errs2 ? 1 : 0;
            err_vec[47] <= (a47 == 8'b0) & errs2 ? 1 : 0;
            err_vec[48] <= (a48 == 8'b0) & errs2 ? 1 : 0;
            err_vec[49] <= (a49 == 8'b0) & errs2 ? 1 : 0;
            err_vec[50] <= (a50 == 8'b0) & errs2 ? 1 : 0;
            err_vec[51] <= (a51 == 8'b0) & errs2 ? 1 : 0;
            err_vec[52] <= (a52 == 8'b0) & errs2 ? 1 : 0;
            err_vec[53] <= (a53 == 8'b0) & errs2 ? 1 : 0;
            err_vec[54] <= (a54 == 8'b0) & errs2 ? 1 : 0;
            err_vec[55] <= (a55 == 8'b0) & errs2 ? 1 : 0;
            err_vec[56] <= (a56 == 8'b0) & errs2 ? 1 : 0;
            err_vec[57] <= (a57 == 8'b0) & errs2 ? 1 : 0;
            err_vec[58] <= (a58 == 8'b0) & errs2 ? 1 : 0;
            err_vec[59] <= (a59 == 8'b0) & errs2 ? 1 : 0;
            err_vec[60] <= (a60 == 8'b0) & errs2 ? 1 : 0;
            err_vec[61] <= (a61 == 8'b0) & errs2 ? 1 : 0;
            err_vec[62] <= (a62 == 8'b0) & errs2 ? 1 : 0;
            err_vec[63] <= (a63 == 8'b0) & errs2 ? 1 : 0;
            err_vec[64] <= (a64 == 8'b0) & errs2 ? 1 : 0;
            err_vec[65] <= (a65 == 8'b0) & errs2 ? 1 : 0;
            err_vec[66] <= (a66 == 8'b0) & errs2 ? 1 : 0;
            err_vec[67] <= (a67 == 8'b0) & errs2 ? 1 : 0;
            err_vec[68] <= (a68 == 8'b0) & errs2 ? 1 : 0;
            err_vec[69] <= (a69 == 8'b0) & errs2 ? 1 : 0;
            err_vec[70] <= (a70 == 8'b0) & errs2 ? 1 : 0;
            err_vec[71] <= (a71 == 8'b0) & errs2 ? 1 : 0;
            err_vec[72] <= (a72 == 8'b0) & errs2 ? 1 : 0;
            err_vec[73] <= (a73 == 8'b0) & errs2 ? 1 : 0;
            err_vec[74] <= (a74 == 8'b0) & errs2 ? 1 : 0;
            err_vec[75] <= (a75 == 8'b0) & errs2 ? 1 : 0;
            err_vec[76] <= (a76 == 8'b0) & errs2 ? 1 : 0;
            err_vec[77] <= (a77 == 8'b0) & errs2 ? 1 : 0;
            err_vec[78] <= (a78 == 8'b0) & errs2 ? 1 : 0;
            err_vec[79] <= (a79 == 8'b0) & errs2 ? 1 : 0;
            err_vec[80] <= (a80 == 8'b0) & errs2 ? 1 : 0;
            err_vec[81] <= (a81 == 8'b0) & errs2 ? 1 : 0;
            err_vec[82] <= (a82 == 8'b0) & errs2 ? 1 : 0;
            err_vec[83] <= (a83 == 8'b0) & errs2 ? 1 : 0;
            err_vec[84] <= (a84 == 8'b0) & errs2 ? 1 : 0;
            err_vec[85] <= (a85 == 8'b0) & errs2 ? 1 : 0;
            err_vec[86] <= (a86 == 8'b0) & errs2 ? 1 : 0;
            err_vec[87] <= (a87 == 8'b0) & errs2 ? 1 : 0;
            err_vec[88] <= (a88 == 8'b0) & errs2 ? 1 : 0;
            err_vec[89] <= (a89 == 8'b0) & errs2 ? 1 : 0;
            err_vec[90] <= (a90 == 8'b0) & errs2 ? 1 : 0;
            err_vec[91] <= (a91 == 8'b0) & errs2 ? 1 : 0;
            err_vec[92] <= (a92 == 8'b0) & errs2 ? 1 : 0;
            err_vec[93] <= (a93 == 8'b0) & errs2 ? 1 : 0;
            err_vec[94] <= (a94 == 8'b0) & errs2 ? 1 : 0;
            err_vec[95] <= (a95 == 8'b0) & errs2 ? 1 : 0;
            err_vec[96] <= (a96 == 8'b0) & errs2 ? 1 : 0;
            err_vec[97] <= (a97 == 8'b0) & errs2 ? 1 : 0;
            err_vec[98] <= (a98 == 8'b0) & errs2 ? 1 : 0;
            err_vec[99] <= (a99 == 8'b0) & errs2 ? 1 : 0;
            err_vec[100] <= (a100 == 8'b0) & errs2 ? 1 : 0;
            err_vec[101] <= (a101 == 8'b0) & errs2 ? 1 : 0;
            err_vec[102] <= (a102 == 8'b0) & errs2 ? 1 : 0;
            err_vec[103] <= (a103 == 8'b0) & errs2 ? 1 : 0;
            err_vec[104] <= (a104 == 8'b0) & errs2 ? 1 : 0;
            err_vec[105] <= (a105 == 8'b0) & errs2 ? 1 : 0;
            err_vec[106] <= (a106 == 8'b0) & errs2 ? 1 : 0;
            err_vec[107] <= (a107 == 8'b0) & errs2 ? 1 : 0;
            err_vec[108] <= (a108 == 8'b0) & errs2 ? 1 : 0;
            err_vec[109] <= (a109 == 8'b0) & errs2 ? 1 : 0;
            err_vec[110] <= (a110 == 8'b0) & errs2 ? 1 : 0;
            err_vec[111] <= (a111 == 8'b0) & errs2 ? 1 : 0;
            err_vec[112] <= (a112 == 8'b0) & errs2 ? 1 : 0;
            err_vec[113] <= (a113 == 8'b0) & errs2 ? 1 : 0;
            err_vec[114] <= (a114 == 8'b0) & errs2 ? 1 : 0;
            err_vec[115] <= (a115 == 8'b0) & errs2 ? 1 : 0;
            err_vec[116] <= (a116 == 8'b0) & errs2 ? 1 : 0;
            err_vec[117] <= (a117 == 8'b0) & errs2 ? 1 : 0;
            err_vec[118] <= (a118 == 8'b0) & errs2 ? 1 : 0;
            err_vec[119] <= (a119 == 8'b0) & errs2 ? 1 : 0;
            err_vec[120] <= (a120 == 8'b0) & errs2 ? 1 : 0;
            err_vec[121] <= (a121 == 8'b0) & errs2 ? 1 : 0;
            err_vec[122] <= (a122 == 8'b0) & errs2 ? 1 : 0;
            err_vec[123] <= (a123 == 8'b0) & errs2 ? 1 : 0;
            err_vec[124] <= (a124 == 8'b0) & errs2 ? 1 : 0;
            err_vec[125] <= (a125 == 8'b0) & errs2 ? 1 : 0;
            err_vec[126] <= (a126 == 8'b0) & errs2 ? 1 : 0;
            err_vec[127] <= (a127 == 8'b0) & errs2 ? 1 : 0;
            err_vec[128] <= (a128 == 8'b0) & errs2 ? 1 : 0;
            err_vec[129] <= (a129 == 8'b0) & errs2 ? 1 : 0;
            err_vec[130] <= (a130 == 8'b0) & errs2 ? 1 : 0;
            err_vec[131] <= (a131 == 8'b0) & errs2 ? 1 : 0;
            err_vec[132] <= (a132 == 8'b0) & errs2 ? 1 : 0;
            err_vec[133] <= (a133 == 8'b0) & errs2 ? 1 : 0;
            err_vec[134] <= (a134 == 8'b0) & errs2 ? 1 : 0;
            err_vec[135] <= (a135 == 8'b0) & errs2 ? 1 : 0;
            err_vec[136] <= (a136 == 8'b0) & errs2 ? 1 : 0;
            err_vec[137] <= (a137 == 8'b0) & errs2 ? 1 : 0;
            err_vec[138] <= (a138 == 8'b0) & errs2 ? 1 : 0;
            err_vec[139] <= (a139 == 8'b0) & errs2 ? 1 : 0;
            err_vec[140] <= (a140 == 8'b0) & errs2 ? 1 : 0;
            err_vec[141] <= (a141 == 8'b0) & errs2 ? 1 : 0;
            err_vec[142] <= (a142 == 8'b0) & errs2 ? 1 : 0;
            err_vec[143] <= (a143 == 8'b0) & errs2 ? 1 : 0;
            err_vec[144] <= (a144 == 8'b0) & errs2 ? 1 : 0;
            err_vec[145] <= (a145 == 8'b0) & errs2 ? 1 : 0;
            err_vec[146] <= (a146 == 8'b0) & errs2 ? 1 : 0;
            err_vec[147] <= (a147 == 8'b0) & errs2 ? 1 : 0;
            err_vec[148] <= (a148 == 8'b0) & errs2 ? 1 : 0;
            err_vec[149] <= (a149 == 8'b0) & errs2 ? 1 : 0;
            err_vec[150] <= (a150 == 8'b0) & errs2 ? 1 : 0;
            err_vec[151] <= (a151 == 8'b0) & errs2 ? 1 : 0;
            err_vec[152] <= (a152 == 8'b0) & errs2 ? 1 : 0;
            err_vec[153] <= (a153 == 8'b0) & errs2 ? 1 : 0;
            err_vec[154] <= (a154 == 8'b0) & errs2 ? 1 : 0;
            err_vec[155] <= (a155 == 8'b0) & errs2 ? 1 : 0;
            err_vec[156] <= (a156 == 8'b0) & errs2 ? 1 : 0;
            err_vec[157] <= (a157 == 8'b0) & errs2 ? 1 : 0;
            err_vec[158] <= (a158 == 8'b0) & errs2 ? 1 : 0;
            err_vec[159] <= (a159 == 8'b0) & errs2 ? 1 : 0;
            err_vec[160] <= (a160 == 8'b0) & errs2 ? 1 : 0;
            err_vec[161] <= (a161 == 8'b0) & errs2 ? 1 : 0;
            err_vec[162] <= (a162 == 8'b0) & errs2 ? 1 : 0;
            err_vec[163] <= (a163 == 8'b0) & errs2 ? 1 : 0;
            err_vec[164] <= (a164 == 8'b0) & errs2 ? 1 : 0;
            err_vec[165] <= (a165 == 8'b0) & errs2 ? 1 : 0;
            err_vec[166] <= (a166 == 8'b0) & errs2 ? 1 : 0;
            err_vec[167] <= (a167 == 8'b0) & errs2 ? 1 : 0;
            err_vec[168] <= (a168 == 8'b0) & errs2 ? 1 : 0;
            err_vec[169] <= (a169 == 8'b0) & errs2 ? 1 : 0;
            err_vec[170] <= (a170 == 8'b0) & errs2 ? 1 : 0;
            err_vec[171] <= (a171 == 8'b0) & errs2 ? 1 : 0;
            err_vec[172] <= (a172 == 8'b0) & errs2 ? 1 : 0;
            err_vec[173] <= (a173 == 8'b0) & errs2 ? 1 : 0;
            err_vec[174] <= (a174 == 8'b0) & errs2 ? 1 : 0;
            err_vec[175] <= (a175 == 8'b0) & errs2 ? 1 : 0;
            err_vec[176] <= (a176 == 8'b0) & errs2 ? 1 : 0;
            err_vec[177] <= (a177 == 8'b0) & errs2 ? 1 : 0;
            err_vec[178] <= (a178 == 8'b0) & errs2 ? 1 : 0;
            err_vec[179] <= (a179 == 8'b0) & errs2 ? 1 : 0;
            err_vec[180] <= (a180 == 8'b0) & errs2 ? 1 : 0;
            err_vec[181] <= (a181 == 8'b0) & errs2 ? 1 : 0;
            err_vec[182] <= (a182 == 8'b0) & errs2 ? 1 : 0;
            err_vec[183] <= (a183 == 8'b0) & errs2 ? 1 : 0;
            err_vec[184] <= (a184 == 8'b0) & errs2 ? 1 : 0;
            err_vec[185] <= (a185 == 8'b0) & errs2 ? 1 : 0;
            err_vec[186] <= (a186 == 8'b0) & errs2 ? 1 : 0;
            err_vec[187] <= (a187 == 8'b0) & errs2 ? 1 : 0;
            err_vec[188] <= (a188 == 8'b0) & errs2 ? 1 : 0;
            err_vec[189] <= (a189 == 8'b0) & errs2 ? 1 : 0;
            err_vec[190] <= (a190 == 8'b0) & errs2 ? 1 : 0;
            err_vec[191] <= (a191 == 8'b0) & errs2 ? 1 : 0;
            err_vec[192] <= (a192 == 8'b0) & errs2 ? 1 : 0;
            err_vec[193] <= (a193 == 8'b0) & errs2 ? 1 : 0;
            err_vec[194] <= (a194 == 8'b0) & errs2 ? 1 : 0;
            err_vec[195] <= (a195 == 8'b0) & errs2 ? 1 : 0;
            err_vec[196] <= (a196 == 8'b0) & errs2 ? 1 : 0;
            err_vec[197] <= (a197 == 8'b0) & errs2 ? 1 : 0;
            err_vec[198] <= (a198 == 8'b0) & errs2 ? 1 : 0;
            err_vec[199] <= (a199 == 8'b0) & errs2 ? 1 : 0;
            err_vec[200] <= (a200 == 8'b0) & errs2 ? 1 : 0;
            err_vec[201] <= (a201 == 8'b0) & errs2 ? 1 : 0;
            err_vec[202] <= (a202 == 8'b0) & errs2 ? 1 : 0;
            err_vec[203] <= (a203 == 8'b0) & errs2 ? 1 : 0;
            err_vec[204] <= (a204 == 8'b0) & errs2 ? 1 : 0;
            err_vec[205] <= (a205 == 8'b0) & errs2 ? 1 : 0;
            err_vec[206] <= (a206 == 8'b0) & errs2 ? 1 : 0;
            err_vec[207] <= (a207 == 8'b0) & errs2 ? 1 : 0;
            err_vec[208] <= (a208 == 8'b0) & errs2 ? 1 : 0;
            err_vec[209] <= (a209 == 8'b0) & errs2 ? 1 : 0;
            err_vec[210] <= (a210 == 8'b0) & errs2 ? 1 : 0;
            err_vec[211] <= (a211 == 8'b0) & errs2 ? 1 : 0;
            err_vec[212] <= (a212 == 8'b0) & errs2 ? 1 : 0;
            err_vec[213] <= (a213 == 8'b0) & errs2 ? 1 : 0;
            err_vec[214] <= (a214 == 8'b0) & errs2 ? 1 : 0;
            err_vec[215] <= (a215 == 8'b0) & errs2 ? 1 : 0;
            err_vec[216] <= (a216 == 8'b0) & errs2 ? 1 : 0;
            err_vec[217] <= (a217 == 8'b0) & errs2 ? 1 : 0;
            err_vec[218] <= (a218 == 8'b0) & errs2 ? 1 : 0;
            err_vec[219] <= (a219 == 8'b0) & errs2 ? 1 : 0;
            err_vec[220] <= (a220 == 8'b0) & errs2 ? 1 : 0;
            err_vec[221] <= (a221 == 8'b0) & errs2 ? 1 : 0;
            err_vec[222] <= (a222 == 8'b0) & errs2 ? 1 : 0;
            err_vec[223] <= (a223 == 8'b0) & errs2 ? 1 : 0;
            err_vec[224] <= (a224 == 8'b0) & errs2 ? 1 : 0;
            err_vec[225] <= (a225 == 8'b0) & errs2 ? 1 : 0;
            err_vec[226] <= (a226 == 8'b0) & errs2 ? 1 : 0;
            err_vec[227] <= (a227 == 8'b0) & errs2 ? 1 : 0;
            err_vec[228] <= (a228 == 8'b0) & errs2 ? 1 : 0;
            err_vec[229] <= (a229 == 8'b0) & errs2 ? 1 : 0;
            err_vec[230] <= (a230 == 8'b0) & errs2 ? 1 : 0;
            err_vec[231] <= (a231 == 8'b0) & errs2 ? 1 : 0;
            err_vec[232] <= (a232 == 8'b0) & errs2 ? 1 : 0;
            err_vec[233] <= (a233 == 8'b0) & errs2 ? 1 : 0;
            err_vec[234] <= (a234 == 8'b0) & errs2 ? 1 : 0;
            err_vec[235] <= (a235 == 8'b0) & errs2 ? 1 : 0;
            err_vec[236] <= (a236 == 8'b0) & errs2 ? 1 : 0;
            err_vec[237] <= (a237 == 8'b0) & errs2 ? 1 : 0;
            err_vec[238] <= (a238 == 8'b0) & errs2 ? 1 : 0;
            err_vec[239] <= (a239 == 8'b0) & errs2 ? 1 : 0;
            err_vec[240] <= (a240 == 8'b0) & errs2 ? 1 : 0;
            err_vec[241] <= (a241 == 8'b0) & errs2 ? 1 : 0;
            err_vec[242] <= (a242 == 8'b0) & errs2 ? 1 : 0;
            err_vec[243] <= (a243 == 8'b0) & errs2 ? 1 : 0;
            err_vec[244] <= (a244 == 8'b0) & errs2 ? 1 : 0;
            err_vec[245] <= (a245 == 8'b0) & errs2 ? 1 : 0;
            err_vec[246] <= (a246 == 8'b0) & errs2 ? 1 : 0;
            err_vec[247] <= (a247 == 8'b0) & errs2 ? 1 : 0;
            err_vec[248] <= (a248 == 8'b0) & errs2 ? 1 : 0;
            err_vec[249] <= (a249 == 8'b0) & errs2 ? 1 : 0;
            err_vec[250] <= (a250 == 8'b0) & errs2 ? 1 : 0;
            err_vec[251] <= (a251 == 8'b0) & errs2 ? 1 : 0;
            err_vec[252] <= (a252 == 8'b0) & errs2 ? 1 : 0;
            err_vec[253] <= (a253 == 8'b0) & errs2 ? 1 : 0;
            err_vec[254] <= (a254 == 8'b0) & errs2 ? 1 : 0;

            
            errs3 <= errs2;
            r4 <= r3;
            
            a0_1  <= a0; 
            a1_1  <= a1; 
            a2_1  <= a2; 
            a3_1  <= a3; 
            a4_1  <= a4; 
            a5_1  <= a5; 
            a6_1  <= a6; 
            a7_1  <= a7; 
            a8_1  <= a8; 
            a9_1  <= a9; 
            a10_1 <= a10; 
            a11_1 <= a11; 
            a12_1 <= a12; 
            a13_1 <= a13; 
            a14_1 <= a14; 
            a15_1 <= a15; 
            a16_1 <= a16; 
            a17_1 <= a17; 
            a18_1 <= a18; 
            a19_1 <= a19; 
            a20_1 <= a20; 
            a21_1 <= a21; 
            a22_1 <= a22; 
            a23_1 <= a23; 
            a24_1 <= a24; 
            a25_1 <= a25; 
            a26_1 <= a26; 
            a27_1 <= a27; 
            a28_1 <= a28; 
            a29_1 <= a29; 
            a30_1 <= a30; 
            a31_1 <= a31; 
            a32_1 <= a32; 
            a33_1 <= a33; 
            a34_1 <= a34; 
            a35_1 <= a35; 
            a36_1 <= a36; 
            a37_1 <= a37; 
            a38_1 <= a38; 
            a39_1 <= a39; 
            a40_1 <= a40; 
            a41_1 <= a41; 
            a42_1 <= a42; 
            a43_1 <= a43; 
            a44_1 <= a44; 
            a45_1 <= a45; 
            a46_1 <= a46; 
            a47_1 <= a47; 
            a48_1 <= a48; 
            a49_1 <= a49; 
            a50_1 <= a50; 
            a51_1 <= a51; 
            a52_1 <= a52; 
            a53_1 <= a53; 
            a54_1 <= a54; 
            a55_1 <= a55; 
            a56_1 <= a56; 
            a57_1 <= a57; 
            a58_1 <= a58; 
            a59_1 <= a59; 
            a60_1 <= a60; 
            a61_1 <= a61; 
            a62_1 <= a62; 
            a63_1 <= a63; 
            a64_1 <= a64; 
            a65_1 <= a65; 
            a66_1 <= a66; 
            a67_1 <= a67; 
            a68_1 <= a68; 
            a69_1 <= a69; 
            a70_1 <= a70; 
            a71_1 <= a71; 
            a72_1 <= a72; 
            a73_1 <= a73; 
            a74_1 <= a74; 
            a75_1 <= a75; 
            a76_1 <= a76; 
            a77_1 <= a77; 
            a78_1 <= a78; 
            a79_1 <= a79; 
            a80_1 <= a80; 
            a81_1 <= a81; 
            a82_1 <= a82; 
            a83_1 <= a83; 
            a84_1 <= a84; 
            a85_1 <= a85; 
            a86_1 <= a86; 
            a87_1 <= a87; 
            a88_1 <= a88; 
            a89_1 <= a89; 
            a90_1 <= a90; 
            a91_1 <= a91; 
            a92_1 <= a92; 
            a93_1 <= a93; 
            a94_1 <= a94; 
            a95_1 <= a95; 
            a96_1 <= a96; 
            a97_1 <= a97; 
            a98_1 <= a98; 
            a99_1 <= a99; 
            a100_1 <= a100; 
            a101_1 <= a101; 
            a102_1 <= a102; 
            a103_1 <= a103; 
            a104_1 <= a104; 
            a105_1 <= a105; 
            a106_1 <= a106; 
            a107_1 <= a107; 
            a108_1 <= a108; 
            a109_1 <= a109; 
            a110_1 <= a110; 
            a111_1 <= a111; 
            a112_1 <= a112; 
            a113_1 <= a113; 
            a114_1 <= a114; 
            a115_1 <= a115; 
            a116_1 <= a116; 
            a117_1 <= a117; 
            a118_1 <= a118; 
            a119_1 <= a119; 
            a120_1 <= a120; 
            a121_1 <= a121; 
            a122_1 <= a122; 
            a123_1 <= a123; 
            a124_1 <= a124; 
            a125_1 <= a125; 
            a126_1 <= a126; 
            a127_1 <= a127; 
            a128_1 <= a128; 
            a129_1 <= a129; 
            a130_1 <= a130; 
            a131_1 <= a131; 
            a132_1 <= a132; 
            a133_1 <= a133; 
            a134_1 <= a134; 
            a135_1 <= a135; 
            a136_1 <= a136; 
            a137_1 <= a137; 
            a138_1 <= a138; 
            a139_1 <= a139; 
            a140_1 <= a140; 
            a141_1 <= a141; 
            a142_1 <= a142; 
            a143_1 <= a143; 
            a144_1 <= a144; 
            a145_1 <= a145; 
            a146_1 <= a146; 
            a147_1 <= a147; 
            a148_1 <= a148; 
            a149_1 <= a149; 
            a150_1 <= a150; 
            a151_1 <= a151; 
            a152_1 <= a152; 
            a153_1 <= a153; 
            a154_1 <= a154; 
            a155_1 <= a155; 
            a156_1 <= a156; 
            a157_1 <= a157; 
            a158_1 <= a158; 
            a159_1 <= a159; 
            a160_1 <= a160; 
            a161_1 <= a161; 
            a162_1 <= a162; 
            a163_1 <= a163; 
            a164_1 <= a164; 
            a165_1 <= a165; 
            a166_1 <= a166; 
            a167_1 <= a167; 
            a168_1 <= a168; 
            a169_1 <= a169; 
            a170_1 <= a170; 
            a171_1 <= a171; 
            a172_1 <= a172; 
            a173_1 <= a173; 
            a174_1 <= a174; 
            a175_1 <= a175; 
            a176_1 <= a176; 
            a177_1 <= a177; 
            a178_1 <= a178; 
            a179_1 <= a179; 
            a180_1 <= a180; 
            a181_1 <= a181; 
            a182_1 <= a182; 
            a183_1 <= a183; 
            a184_1 <= a184; 
            a185_1 <= a185; 
            a186_1 <= a186; 
            a187_1 <= a187; 
            a188_1 <= a188; 
            a189_1 <= a189; 
            a190_1 <= a190; 
            a191_1 <= a191; 
            a192_1 <= a192; 
            a193_1 <= a193; 
            a194_1 <= a194; 
            a195_1 <= a195; 
            a196_1 <= a196; 
            a197_1 <= a197; 
            a198_1 <= a198; 
            a199_1 <= a199; 
            a200_1 <= a200; 
            a201_1 <= a201; 
            a202_1 <= a202; 
            a203_1 <= a203; 
            a204_1 <= a204; 
            a205_1 <= a205; 
            a206_1 <= a206; 
            a207_1 <= a207; 
            a208_1 <= a208; 
            a209_1 <= a209; 
            a210_1 <= a210; 
            a211_1 <= a211; 
            a212_1 <= a212; 
            a213_1 <= a213; 
            a214_1 <= a214; 
            a215_1 <= a215; 
            a216_1 <= a216; 
            a217_1 <= a217; 
            a218_1 <= a218; 
            a219_1 <= a219; 
            a220_1 <= a220; 
            a221_1 <= a221; 
            a222_1 <= a222; 
            a223_1 <= a223; 
            a224_1 <= a224; 
            a225_1 <= a225; 
            a226_1 <= a226; 
            a227_1 <= a227; 
            a228_1 <= a228; 
            a229_1 <= a229; 
            a230_1 <= a230; 
            a231_1 <= a231; 
            a232_1 <= a232; 
            a233_1 <= a233; 
            a234_1 <= a234; 
            a235_1 <= a235; 
            a236_1 <= a236; 
            a237_1 <= a237; 
            a238_1 <= a238; 
            a239_1 <= a239; 
            a240_1 <= a240; 
            a241_1 <= a241; 
            a242_1 <= a242; 
            a243_1 <= a243; 
            a244_1 <= a244; 
            a245_1 <= a245; 
            a246_1 <= a246; 
            a247_1 <= a247; 
            a248_1 <= a248; 
            a249_1 <= a249; 
            a250_1 <= a250; 
            a251_1 <= a251; 
            a252_1 <= a252; 
            a253_1 <= a253; 
            a254_1 <= a254; 

            
            //Clock Cycle 5: Count errors
            for (x=0,temp=0; x<255; x=x+1) begin
                temp = temp + err_vec[x];
            end

            d <= temp;
            d_e <= (temp + (^r4)) % 2;
            
            errs4 <= errs3;
            r5 <= r4;
            
            a0_2 <= a0_1; 
            a1_2 <= a1_1; 
            a2_2 <= a2_1; 
            a3_2 <= a3_1; 
            a4_2 <= a4_1; 
            a5_2 <= a5_1; 
            a6_2 <= a6_1; 
            a7_2 <= a7_1; 
            a8_2 <= a8_1; 
            a9_2 <= a9_1; 
            a10_2 <= a10_1; 
            a11_2 <= a11_1; 
            a12_2 <= a12_1; 
            a13_2 <= a13_1; 
            a14_2 <= a14_1; 
            a15_2 <= a15_1; 
            a16_2 <= a16_1; 
            a17_2 <= a17_1; 
            a18_2 <= a18_1; 
            a19_2 <= a19_1; 
            a20_2 <= a20_1; 
            a21_2 <= a21_1; 
            a22_2 <= a22_1; 
            a23_2 <= a23_1; 
            a24_2 <= a24_1; 
            a25_2 <= a25_1; 
            a26_2 <= a26_1; 
            a27_2 <= a27_1; 
            a28_2 <= a28_1; 
            a29_2 <= a29_1; 
            a30_2 <= a30_1; 
            a31_2 <= a31_1; 
            a32_2 <= a32_1; 
            a33_2 <= a33_1; 
            a34_2 <= a34_1; 
            a35_2 <= a35_1; 
            a36_2 <= a36_1; 
            a37_2 <= a37_1; 
            a38_2 <= a38_1; 
            a39_2 <= a39_1; 
            a40_2 <= a40_1; 
            a41_2 <= a41_1; 
            a42_2 <= a42_1; 
            a43_2 <= a43_1; 
            a44_2 <= a44_1; 
            a45_2 <= a45_1; 
            a46_2 <= a46_1; 
            a47_2 <= a47_1; 
            a48_2 <= a48_1; 
            a49_2 <= a49_1; 
            a50_2 <= a50_1; 
            a51_2 <= a51_1; 
            a52_2 <= a52_1; 
            a53_2 <= a53_1; 
            a54_2 <= a54_1; 
            a55_2 <= a55_1; 
            a56_2 <= a56_1; 
            a57_2 <= a57_1; 
            a58_2 <= a58_1; 
            a59_2 <= a59_1; 
            a60_2 <= a60_1; 
            a61_2 <= a61_1; 
            a62_2 <= a62_1; 
            a63_2 <= a63_1; 
            a64_2 <= a64_1; 
            a65_2 <= a65_1; 
            a66_2 <= a66_1; 
            a67_2 <= a67_1; 
            a68_2 <= a68_1; 
            a69_2 <= a69_1; 
            a70_2 <= a70_1; 
            a71_2 <= a71_1; 
            a72_2 <= a72_1; 
            a73_2 <= a73_1; 
            a74_2 <= a74_1; 
            a75_2 <= a75_1; 
            a76_2 <= a76_1; 
            a77_2 <= a77_1; 
            a78_2 <= a78_1; 
            a79_2 <= a79_1; 
            a80_2 <= a80_1; 
            a81_2 <= a81_1; 
            a82_2 <= a82_1; 
            a83_2 <= a83_1; 
            a84_2 <= a84_1; 
            a85_2 <= a85_1; 
            a86_2 <= a86_1; 
            a87_2 <= a87_1; 
            a88_2 <= a88_1; 
            a89_2 <= a89_1; 
            a90_2 <= a90_1; 
            a91_2 <= a91_1; 
            a92_2 <= a92_1; 
            a93_2 <= a93_1; 
            a94_2 <= a94_1; 
            a95_2 <= a95_1; 
            a96_2 <= a96_1; 
            a97_2 <= a97_1; 
            a98_2 <= a98_1; 
            a99_2 <= a99_1; 
            a100_2 <= a100_1; 
            a101_2 <= a101_1; 
            a102_2 <= a102_1; 
            a103_2 <= a103_1; 
            a104_2 <= a104_1; 
            a105_2 <= a105_1; 
            a106_2 <= a106_1; 
            a107_2 <= a107_1; 
            a108_2 <= a108_1; 
            a109_2 <= a109_1; 
            a110_2 <= a110_1; 
            a111_2 <= a111_1; 
            a112_2 <= a112_1; 
            a113_2 <= a113_1; 
            a114_2 <= a114_1; 
            a115_2 <= a115_1; 
            a116_2 <= a116_1; 
            a117_2 <= a117_1; 
            a118_2 <= a118_1; 
            a119_2 <= a119_1; 
            a120_2 <= a120_1; 
            a121_2 <= a121_1; 
            a122_2 <= a122_1; 
            a123_2 <= a123_1; 
            a124_2 <= a124_1; 
            a125_2 <= a125_1; 
            a126_2 <= a126_1; 
            a127_2 <= a127_1; 
            a128_2 <= a128_1; 
            a129_2 <= a129_1; 
            a130_2 <= a130_1; 
            a131_2 <= a131_1; 
            a132_2 <= a132_1; 
            a133_2 <= a133_1; 
            a134_2 <= a134_1; 
            a135_2 <= a135_1; 
            a136_2 <= a136_1; 
            a137_2 <= a137_1; 
            a138_2 <= a138_1; 
            a139_2 <= a139_1; 
            a140_2 <= a140_1; 
            a141_2 <= a141_1; 
            a142_2 <= a142_1; 
            a143_2 <= a143_1; 
            a144_2 <= a144_1; 
            a145_2 <= a145_1; 
            a146_2 <= a146_1; 
            a147_2 <= a147_1; 
            a148_2 <= a148_1; 
            a149_2 <= a149_1; 
            a150_2 <= a150_1; 
            a151_2 <= a151_1; 
            a152_2 <= a152_1; 
            a153_2 <= a153_1; 
            a154_2 <= a154_1; 
            a155_2 <= a155_1; 
            a156_2 <= a156_1; 
            a157_2 <= a157_1; 
            a158_2 <= a158_1; 
            a159_2 <= a159_1; 
            a160_2 <= a160_1; 
            a161_2 <= a161_1; 
            a162_2 <= a162_1; 
            a163_2 <= a163_1; 
            a164_2 <= a164_1; 
            a165_2 <= a165_1; 
            a166_2 <= a166_1; 
            a167_2 <= a167_1; 
            a168_2 <= a168_1; 
            a169_2 <= a169_1; 
            a170_2 <= a170_1; 
            a171_2 <= a171_1; 
            a172_2 <= a172_1; 
            a173_2 <= a173_1; 
            a174_2 <= a174_1; 
            a175_2 <= a175_1; 
            a176_2 <= a176_1; 
            a177_2 <= a177_1; 
            a178_2 <= a178_1; 
            a179_2 <= a179_1; 
            a180_2 <= a180_1; 
            a181_2 <= a181_1; 
            a182_2 <= a182_1; 
            a183_2 <= a183_1; 
            a184_2 <= a184_1; 
            a185_2 <= a185_1; 
            a186_2 <= a186_1; 
            a187_2 <= a187_1; 
            a188_2 <= a188_1; 
            a189_2 <= a189_1; 
            a190_2 <= a190_1; 
            a191_2 <= a191_1; 
            a192_2 <= a192_1; 
            a193_2 <= a193_1; 
            a194_2 <= a194_1; 
            a195_2 <= a195_1; 
            a196_2 <= a196_1; 
            a197_2 <= a197_1; 
            a198_2 <= a198_1; 
            a199_2 <= a199_1; 
            a200_2 <= a200_1; 
            a201_2 <= a201_1; 
            a202_2 <= a202_1; 
            a203_2 <= a203_1; 
            a204_2 <= a204_1; 
            a205_2 <= a205_1; 
            a206_2 <= a206_1; 
            a207_2 <= a207_1; 
            a208_2 <= a208_1; 
            a209_2 <= a209_1; 
            a210_2 <= a210_1; 
            a211_2 <= a211_1; 
            a212_2 <= a212_1; 
            a213_2 <= a213_1; 
            a214_2 <= a214_1; 
            a215_2 <= a215_1; 
            a216_2 <= a216_1; 
            a217_2 <= a217_1; 
            a218_2 <= a218_1; 
            a219_2 <= a219_1; 
            a220_2 <= a220_1; 
            a221_2 <= a221_1; 
            a222_2 <= a222_1; 
            a223_2 <= a223_1; 
            a224_2 <= a224_1; 
            a225_2 <= a225_1; 
            a226_2 <= a226_1; 
            a227_2 <= a227_1; 
            a228_2 <= a228_1; 
            a229_2 <= a229_1; 
            a230_2 <= a230_1; 
            a231_2 <= a231_1; 
            a232_2 <= a232_1; 
            a233_2 <= a233_1; 
            a234_2 <= a234_1; 
            a235_2 <= a235_1; 
            a236_2 <= a236_1; 
            a237_2 <= a237_1; 
            a238_2 <= a238_1; 
            a239_2 <= a239_1; 
            a240_2 <= a240_1; 
            a241_2 <= a241_1; 
            a242_2 <= a242_1; 
            a243_2 <= a243_1; 
            a244_2 <= a244_1; 
            a245_2 <= a245_1; 
            a246_2 <= a246_1; 
            a247_2 <= a247_1; 
            a248_2 <= a248_1; 
            a249_2 <= a249_1; 
            a250_2 <= a250_1; 
            a251_2 <= a251_1; 
            a252_2 <= a252_1; 
            a253_2 <= a253_1; 
            a254_2 <= a254_1; 

            
            //Clock Cycle 6: Correct errors
//            if(!(d & d_e)) begin
            if (d + d_e <= 2) begin
            
                dec[0]  <= (a0_2  == 8'b0) & errs4 ? ~r5[0] : r5[0]; 
                dec[1]  <= (a1_2  == 8'b0) & errs4 ? ~r5[1] : r5[1]; 
                dec[2]  <= (a2_2  == 8'b0) & errs4 ? ~r5[2] : r5[2]; 
                dec[3]  <= (a3_2  == 8'b0) & errs4 ? ~r5[3] : r5[3]; 
                dec[4]  <= (a4_2  == 8'b0) & errs4 ? ~r5[4] : r5[4]; 
                dec[5]  <= (a5_2  == 8'b0) & errs4 ? ~r5[5] : r5[5]; 
                dec[6]  <= (a6_2  == 8'b0) & errs4 ? ~r5[6] : r5[6]; 
                dec[7]  <= (a7_2  == 8'b0) & errs4 ? ~r5[7] : r5[7]; 
                dec[8]  <= (a8_2  == 8'b0) & errs4 ? ~r5[8] : r5[8]; 
                dec[9]  <= (a9_2  == 8'b0) & errs4 ? ~r5[9] : r5[9]; 
                dec[10] <= (a10_2 == 8'b0) & errs4 ? ~r5[10] : r5[10]; 
                dec[11] <= (a11_2 == 8'b0) & errs4 ? ~r5[11] : r5[11]; 
                dec[12] <= (a12_2 == 8'b0) & errs4 ? ~r5[12] : r5[12]; 
                dec[13] <= (a13_2 == 8'b0) & errs4 ? ~r5[13] : r5[13]; 
                dec[14] <= (a14_2 == 8'b0) & errs4 ? ~r5[14] : r5[14]; 
                dec[15] <= (a15_2 == 8'b0) & errs4 ? ~r5[15] : r5[15]; 
                dec[16] <= (a16_2 == 8'b0) & errs4 ? ~r5[16] : r5[16]; 
                dec[17] <= (a17_2 == 8'b0) & errs4 ? ~r5[17] : r5[17]; 
                dec[18] <= (a18_2 == 8'b0) & errs4 ? ~r5[18] : r5[18]; 
                dec[19] <= (a19_2 == 8'b0) & errs4 ? ~r5[19] : r5[19]; 
                dec[20] <= (a20_2 == 8'b0) & errs4 ? ~r5[20] : r5[20]; 
                dec[21] <= (a21_2 == 8'b0) & errs4 ? ~r5[21] : r5[21]; 
                dec[22] <= (a22_2 == 8'b0) & errs4 ? ~r5[22] : r5[22]; 
                dec[23] <= (a23_2 == 8'b0) & errs4 ? ~r5[23] : r5[23]; 
                dec[24] <= (a24_2 == 8'b0) & errs4 ? ~r5[24] : r5[24]; 
                dec[25] <= (a25_2 == 8'b0) & errs4 ? ~r5[25] : r5[25]; 
                dec[26] <= (a26_2 == 8'b0) & errs4 ? ~r5[26] : r5[26]; 
                dec[27] <= (a27_2 == 8'b0) & errs4 ? ~r5[27] : r5[27]; 
                dec[28] <= (a28_2 == 8'b0) & errs4 ? ~r5[28] : r5[28]; 
                dec[29] <= (a29_2 == 8'b0) & errs4 ? ~r5[29] : r5[29]; 
                dec[30] <= (a30_2 == 8'b0) & errs4 ? ~r5[30] : r5[30]; 
                dec[31] <= (a31_2 == 8'b0) & errs4 ? ~r5[31] : r5[31]; 
                dec[32] <= (a32_2 == 8'b0) & errs4 ? ~r5[32] : r5[32]; 
                dec[33] <= (a33_2 == 8'b0) & errs4 ? ~r5[33] : r5[33]; 
                dec[34] <= (a34_2 == 8'b0) & errs4 ? ~r5[34] : r5[34]; 
                dec[35] <= (a35_2 == 8'b0) & errs4 ? ~r5[35] : r5[35]; 
                dec[36] <= (a36_2 == 8'b0) & errs4 ? ~r5[36] : r5[36]; 
                dec[37] <= (a37_2 == 8'b0) & errs4 ? ~r5[37] : r5[37]; 
                dec[38] <= (a38_2 == 8'b0) & errs4 ? ~r5[38] : r5[38]; 
                dec[39] <= (a39_2 == 8'b0) & errs4 ? ~r5[39] : r5[39]; 
                dec[40] <= (a40_2 == 8'b0) & errs4 ? ~r5[40] : r5[40]; 
                dec[41] <= (a41_2 == 8'b0) & errs4 ? ~r5[41] : r5[41]; 
                dec[42] <= (a42_2 == 8'b0) & errs4 ? ~r5[42] : r5[42]; 
                dec[43] <= (a43_2 == 8'b0) & errs4 ? ~r5[43] : r5[43]; 
                dec[44] <= (a44_2 == 8'b0) & errs4 ? ~r5[44] : r5[44]; 
                dec[45] <= (a45_2 == 8'b0) & errs4 ? ~r5[45] : r5[45]; 
                dec[46] <= (a46_2 == 8'b0) & errs4 ? ~r5[46] : r5[46]; 
                dec[47] <= (a47_2 == 8'b0) & errs4 ? ~r5[47] : r5[47]; 
                dec[48] <= (a48_2 == 8'b0) & errs4 ? ~r5[48] : r5[48]; 
                dec[49] <= (a49_2 == 8'b0) & errs4 ? ~r5[49] : r5[49]; 
                dec[50] <= (a50_2 == 8'b0) & errs4 ? ~r5[50] : r5[50]; 
                dec[51] <= (a51_2 == 8'b0) & errs4 ? ~r5[51] : r5[51]; 
                dec[52] <= (a52_2 == 8'b0) & errs4 ? ~r5[52] : r5[52]; 
                dec[53] <= (a53_2 == 8'b0) & errs4 ? ~r5[53] : r5[53]; 
                dec[54] <= (a54_2 == 8'b0) & errs4 ? ~r5[54] : r5[54]; 
                dec[55] <= (a55_2 == 8'b0) & errs4 ? ~r5[55] : r5[55]; 
                dec[56] <= (a56_2 == 8'b0) & errs4 ? ~r5[56] : r5[56]; 
                dec[57] <= (a57_2 == 8'b0) & errs4 ? ~r5[57] : r5[57]; 
                dec[58] <= (a58_2 == 8'b0) & errs4 ? ~r5[58] : r5[58]; 
                dec[59] <= (a59_2 == 8'b0) & errs4 ? ~r5[59] : r5[59]; 
                dec[60] <= (a60_2 == 8'b0) & errs4 ? ~r5[60] : r5[60]; 
                dec[61] <= (a61_2 == 8'b0) & errs4 ? ~r5[61] : r5[61]; 
                dec[62] <= (a62_2 == 8'b0) & errs4 ? ~r5[62] : r5[62]; 
                dec[63] <= (a63_2 == 8'b0) & errs4 ? ~r5[63] : r5[63]; 
                dec[64] <= (a64_2 == 8'b0) & errs4 ? ~r5[64] : r5[64]; 
                dec[65] <= (a65_2 == 8'b0) & errs4 ? ~r5[65] : r5[65]; 
                dec[66] <= (a66_2 == 8'b0) & errs4 ? ~r5[66] : r5[66]; 
                dec[67] <= (a67_2 == 8'b0) & errs4 ? ~r5[67] : r5[67]; 
                dec[68] <= (a68_2 == 8'b0) & errs4 ? ~r5[68] : r5[68]; 
                dec[69] <= (a69_2 == 8'b0) & errs4 ? ~r5[69] : r5[69]; 
                dec[70] <= (a70_2 == 8'b0) & errs4 ? ~r5[70] : r5[70]; 
                dec[71] <= (a71_2 == 8'b0) & errs4 ? ~r5[71] : r5[71]; 
                dec[72] <= (a72_2 == 8'b0) & errs4 ? ~r5[72] : r5[72]; 
                dec[73] <= (a73_2 == 8'b0) & errs4 ? ~r5[73] : r5[73]; 
                dec[74] <= (a74_2 == 8'b0) & errs4 ? ~r5[74] : r5[74]; 
                dec[75] <= (a75_2 == 8'b0) & errs4 ? ~r5[75] : r5[75]; 
                dec[76] <= (a76_2 == 8'b0) & errs4 ? ~r5[76] : r5[76]; 
                dec[77] <= (a77_2 == 8'b0) & errs4 ? ~r5[77] : r5[77]; 
                dec[78] <= (a78_2 == 8'b0) & errs4 ? ~r5[78] : r5[78]; 
                dec[79] <= (a79_2 == 8'b0) & errs4 ? ~r5[79] : r5[79]; 
                dec[80] <= (a80_2 == 8'b0) & errs4 ? ~r5[80] : r5[80]; 
                dec[81] <= (a81_2 == 8'b0) & errs4 ? ~r5[81] : r5[81]; 
                dec[82] <= (a82_2 == 8'b0) & errs4 ? ~r5[82] : r5[82]; 
                dec[83] <= (a83_2 == 8'b0) & errs4 ? ~r5[83] : r5[83]; 
                dec[84] <= (a84_2 == 8'b0) & errs4 ? ~r5[84] : r5[84]; 
                dec[85] <= (a85_2 == 8'b0) & errs4 ? ~r5[85] : r5[85]; 
                dec[86] <= (a86_2 == 8'b0) & errs4 ? ~r5[86] : r5[86]; 
                dec[87] <= (a87_2 == 8'b0) & errs4 ? ~r5[87] : r5[87]; 
                dec[88] <= (a88_2 == 8'b0) & errs4 ? ~r5[88] : r5[88]; 
                dec[89] <= (a89_2 == 8'b0) & errs4 ? ~r5[89] : r5[89]; 
                dec[90] <= (a90_2 == 8'b0) & errs4 ? ~r5[90] : r5[90]; 
                dec[91] <= (a91_2 == 8'b0) & errs4 ? ~r5[91] : r5[91]; 
                dec[92] <= (a92_2 == 8'b0) & errs4 ? ~r5[92] : r5[92]; 
                dec[93] <= (a93_2 == 8'b0) & errs4 ? ~r5[93] : r5[93]; 
                dec[94] <= (a94_2 == 8'b0) & errs4 ? ~r5[94] : r5[94]; 
                dec[95] <= (a95_2 == 8'b0) & errs4 ? ~r5[95] : r5[95]; 
                dec[96] <= (a96_2 == 8'b0) & errs4 ? ~r5[96] : r5[96]; 
                dec[97] <= (a97_2 == 8'b0) & errs4 ? ~r5[97] : r5[97]; 
                dec[98] <= (a98_2 == 8'b0) & errs4 ? ~r5[98] : r5[98]; 
                dec[99] <= (a99_2 == 8'b0) & errs4 ? ~r5[99] : r5[99]; 
                dec[100] <= (a100_2 == 8'b0) & errs4 ? ~r5[100] : r5[100]; 
                dec[101] <= (a101_2 == 8'b0) & errs4 ? ~r5[101] : r5[101]; 
                dec[102] <= (a102_2 == 8'b0) & errs4 ? ~r5[102] : r5[102]; 
                dec[103] <= (a103_2 == 8'b0) & errs4 ? ~r5[103] : r5[103]; 
                dec[104] <= (a104_2 == 8'b0) & errs4 ? ~r5[104] : r5[104]; 
                dec[105] <= (a105_2 == 8'b0) & errs4 ? ~r5[105] : r5[105]; 
                dec[106] <= (a106_2 == 8'b0) & errs4 ? ~r5[106] : r5[106]; 
                dec[107] <= (a107_2 == 8'b0) & errs4 ? ~r5[107] : r5[107]; 
                dec[108] <= (a108_2 == 8'b0) & errs4 ? ~r5[108] : r5[108]; 
                dec[109] <= (a109_2 == 8'b0) & errs4 ? ~r5[109] : r5[109]; 
                dec[110] <= (a110_2 == 8'b0) & errs4 ? ~r5[110] : r5[110]; 
                dec[111] <= (a111_2 == 8'b0) & errs4 ? ~r5[111] : r5[111]; 
                dec[112] <= (a112_2 == 8'b0) & errs4 ? ~r5[112] : r5[112]; 
                dec[113] <= (a113_2 == 8'b0) & errs4 ? ~r5[113] : r5[113]; 
                dec[114] <= (a114_2 == 8'b0) & errs4 ? ~r5[114] : r5[114]; 
                dec[115] <= (a115_2 == 8'b0) & errs4 ? ~r5[115] : r5[115]; 
                dec[116] <= (a116_2 == 8'b0) & errs4 ? ~r5[116] : r5[116]; 
                dec[117] <= (a117_2 == 8'b0) & errs4 ? ~r5[117] : r5[117]; 
                dec[118] <= (a118_2 == 8'b0) & errs4 ? ~r5[118] : r5[118]; 
                dec[119] <= (a119_2 == 8'b0) & errs4 ? ~r5[119] : r5[119]; 
                dec[120] <= (a120_2 == 8'b0) & errs4 ? ~r5[120] : r5[120]; 
                dec[121] <= (a121_2 == 8'b0) & errs4 ? ~r5[121] : r5[121]; 
                dec[122] <= (a122_2 == 8'b0) & errs4 ? ~r5[122] : r5[122]; 
                dec[123] <= (a123_2 == 8'b0) & errs4 ? ~r5[123] : r5[123]; 
                dec[124] <= (a124_2 == 8'b0) & errs4 ? ~r5[124] : r5[124]; 
                dec[125] <= (a125_2 == 8'b0) & errs4 ? ~r5[125] : r5[125]; 
                dec[126] <= (a126_2 == 8'b0) & errs4 ? ~r5[126] : r5[126]; 
                dec[127] <= (a127_2 == 8'b0) & errs4 ? ~r5[127] : r5[127]; 
                dec[128] <= (a128_2 == 8'b0) & errs4 ? ~r5[128] : r5[128]; 
                dec[129] <= (a129_2 == 8'b0) & errs4 ? ~r5[129] : r5[129]; 
                dec[130] <= (a130_2 == 8'b0) & errs4 ? ~r5[130] : r5[130]; 
                dec[131] <= (a131_2 == 8'b0) & errs4 ? ~r5[131] : r5[131]; 
                dec[132] <= (a132_2 == 8'b0) & errs4 ? ~r5[132] : r5[132]; 
                dec[133] <= (a133_2 == 8'b0) & errs4 ? ~r5[133] : r5[133]; 
                dec[134] <= (a134_2 == 8'b0) & errs4 ? ~r5[134] : r5[134]; 
                dec[135] <= (a135_2 == 8'b0) & errs4 ? ~r5[135] : r5[135]; 
                dec[136] <= (a136_2 == 8'b0) & errs4 ? ~r5[136] : r5[136]; 
                dec[137] <= (a137_2 == 8'b0) & errs4 ? ~r5[137] : r5[137]; 
                dec[138] <= (a138_2 == 8'b0) & errs4 ? ~r5[138] : r5[138]; 
                dec[139] <= (a139_2 == 8'b0) & errs4 ? ~r5[139] : r5[139]; 
                dec[140] <= (a140_2 == 8'b0) & errs4 ? ~r5[140] : r5[140]; 
                dec[141] <= (a141_2 == 8'b0) & errs4 ? ~r5[141] : r5[141]; 
                dec[142] <= (a142_2 == 8'b0) & errs4 ? ~r5[142] : r5[142]; 
                dec[143] <= (a143_2 == 8'b0) & errs4 ? ~r5[143] : r5[143]; 
                dec[144] <= (a144_2 == 8'b0) & errs4 ? ~r5[144] : r5[144]; 
                dec[145] <= (a145_2 == 8'b0) & errs4 ? ~r5[145] : r5[145]; 
                dec[146] <= (a146_2 == 8'b0) & errs4 ? ~r5[146] : r5[146]; 
                dec[147] <= (a147_2 == 8'b0) & errs4 ? ~r5[147] : r5[147]; 
                dec[148] <= (a148_2 == 8'b0) & errs4 ? ~r5[148] : r5[148]; 
                dec[149] <= (a149_2 == 8'b0) & errs4 ? ~r5[149] : r5[149]; 
                dec[150] <= (a150_2 == 8'b0) & errs4 ? ~r5[150] : r5[150]; 
                dec[151] <= (a151_2 == 8'b0) & errs4 ? ~r5[151] : r5[151]; 
                dec[152] <= (a152_2 == 8'b0) & errs4 ? ~r5[152] : r5[152]; 
                dec[153] <= (a153_2 == 8'b0) & errs4 ? ~r5[153] : r5[153]; 
                dec[154] <= (a154_2 == 8'b0) & errs4 ? ~r5[154] : r5[154]; 
                dec[155] <= (a155_2 == 8'b0) & errs4 ? ~r5[155] : r5[155]; 
                dec[156] <= (a156_2 == 8'b0) & errs4 ? ~r5[156] : r5[156]; 
                dec[157] <= (a157_2 == 8'b0) & errs4 ? ~r5[157] : r5[157]; 
                dec[158] <= (a158_2 == 8'b0) & errs4 ? ~r5[158] : r5[158]; 
                dec[159] <= (a159_2 == 8'b0) & errs4 ? ~r5[159] : r5[159]; 
                dec[160] <= (a160_2 == 8'b0) & errs4 ? ~r5[160] : r5[160]; 
                dec[161] <= (a161_2 == 8'b0) & errs4 ? ~r5[161] : r5[161]; 
                dec[162] <= (a162_2 == 8'b0) & errs4 ? ~r5[162] : r5[162]; 
                dec[163] <= (a163_2 == 8'b0) & errs4 ? ~r5[163] : r5[163]; 
                dec[164] <= (a164_2 == 8'b0) & errs4 ? ~r5[164] : r5[164]; 
                dec[165] <= (a165_2 == 8'b0) & errs4 ? ~r5[165] : r5[165]; 
                dec[166] <= (a166_2 == 8'b0) & errs4 ? ~r5[166] : r5[166]; 
                dec[167] <= (a167_2 == 8'b0) & errs4 ? ~r5[167] : r5[167]; 
                dec[168] <= (a168_2 == 8'b0) & errs4 ? ~r5[168] : r5[168]; 
                dec[169] <= (a169_2 == 8'b0) & errs4 ? ~r5[169] : r5[169]; 
                dec[170] <= (a170_2 == 8'b0) & errs4 ? ~r5[170] : r5[170]; 
                dec[171] <= (a171_2 == 8'b0) & errs4 ? ~r5[171] : r5[171]; 
                dec[172] <= (a172_2 == 8'b0) & errs4 ? ~r5[172] : r5[172]; 
                dec[173] <= (a173_2 == 8'b0) & errs4 ? ~r5[173] : r5[173]; 
                dec[174] <= (a174_2 == 8'b0) & errs4 ? ~r5[174] : r5[174]; 
                dec[175] <= (a175_2 == 8'b0) & errs4 ? ~r5[175] : r5[175]; 
                dec[176] <= (a176_2 == 8'b0) & errs4 ? ~r5[176] : r5[176]; 
                dec[177] <= (a177_2 == 8'b0) & errs4 ? ~r5[177] : r5[177]; 
                dec[178] <= (a178_2 == 8'b0) & errs4 ? ~r5[178] : r5[178]; 
                dec[179] <= (a179_2 == 8'b0) & errs4 ? ~r5[179] : r5[179]; 
                dec[180] <= (a180_2 == 8'b0) & errs4 ? ~r5[180] : r5[180]; 
                dec[181] <= (a181_2 == 8'b0) & errs4 ? ~r5[181] : r5[181]; 
                dec[182] <= (a182_2 == 8'b0) & errs4 ? ~r5[182] : r5[182]; 
                dec[183] <= (a183_2 == 8'b0) & errs4 ? ~r5[183] : r5[183]; 
                dec[184] <= (a184_2 == 8'b0) & errs4 ? ~r5[184] : r5[184]; 
                dec[185] <= (a185_2 == 8'b0) & errs4 ? ~r5[185] : r5[185]; 
                dec[186] <= (a186_2 == 8'b0) & errs4 ? ~r5[186] : r5[186]; 
                dec[187] <= (a187_2 == 8'b0) & errs4 ? ~r5[187] : r5[187]; 
                dec[188] <= (a188_2 == 8'b0) & errs4 ? ~r5[188] : r5[188]; 
                dec[189] <= (a189_2 == 8'b0) & errs4 ? ~r5[189] : r5[189]; 
                dec[190] <= (a190_2 == 8'b0) & errs4 ? ~r5[190] : r5[190]; 
                dec[191] <= (a191_2 == 8'b0) & errs4 ? ~r5[191] : r5[191]; 
                dec[192] <= (a192_2 == 8'b0) & errs4 ? ~r5[192] : r5[192]; 
                dec[193] <= (a193_2 == 8'b0) & errs4 ? ~r5[193] : r5[193]; 
                dec[194] <= (a194_2 == 8'b0) & errs4 ? ~r5[194] : r5[194]; 
                dec[195] <= (a195_2 == 8'b0) & errs4 ? ~r5[195] : r5[195]; 
                dec[196] <= (a196_2 == 8'b0) & errs4 ? ~r5[196] : r5[196]; 
                dec[197] <= (a197_2 == 8'b0) & errs4 ? ~r5[197] : r5[197]; 
                dec[198] <= (a198_2 == 8'b0) & errs4 ? ~r5[198] : r5[198]; 
                dec[199] <= (a199_2 == 8'b0) & errs4 ? ~r5[199] : r5[199]; 
                dec[200] <= (a200_2 == 8'b0) & errs4 ? ~r5[200] : r5[200]; 
                dec[201] <= (a201_2 == 8'b0) & errs4 ? ~r5[201] : r5[201]; 
                dec[202] <= (a202_2 == 8'b0) & errs4 ? ~r5[202] : r5[202]; 
                dec[203] <= (a203_2 == 8'b0) & errs4 ? ~r5[203] : r5[203]; 
                dec[204] <= (a204_2 == 8'b0) & errs4 ? ~r5[204] : r5[204]; 
                dec[205] <= (a205_2 == 8'b0) & errs4 ? ~r5[205] : r5[205]; 
                dec[206] <= (a206_2 == 8'b0) & errs4 ? ~r5[206] : r5[206]; 
                dec[207] <= (a207_2 == 8'b0) & errs4 ? ~r5[207] : r5[207]; 
                dec[208] <= (a208_2 == 8'b0) & errs4 ? ~r5[208] : r5[208]; 
                dec[209] <= (a209_2 == 8'b0) & errs4 ? ~r5[209] : r5[209]; 
                dec[210] <= (a210_2 == 8'b0) & errs4 ? ~r5[210] : r5[210]; 
                dec[211] <= (a211_2 == 8'b0) & errs4 ? ~r5[211] : r5[211]; 
                dec[212] <= (a212_2 == 8'b0) & errs4 ? ~r5[212] : r5[212]; 
                dec[213] <= (a213_2 == 8'b0) & errs4 ? ~r5[213] : r5[213]; 
                dec[214] <= (a214_2 == 8'b0) & errs4 ? ~r5[214] : r5[214]; 
                dec[215] <= (a215_2 == 8'b0) & errs4 ? ~r5[215] : r5[215]; 
                dec[216] <= (a216_2 == 8'b0) & errs4 ? ~r5[216] : r5[216]; 
                dec[217] <= (a217_2 == 8'b0) & errs4 ? ~r5[217] : r5[217]; 
                dec[218] <= (a218_2 == 8'b0) & errs4 ? ~r5[218] : r5[218]; 
                dec[219] <= (a219_2 == 8'b0) & errs4 ? ~r5[219] : r5[219]; 
                dec[220] <= (a220_2 == 8'b0) & errs4 ? ~r5[220] : r5[220]; 
                dec[221] <= (a221_2 == 8'b0) & errs4 ? ~r5[221] : r5[221]; 
                dec[222] <= (a222_2 == 8'b0) & errs4 ? ~r5[222] : r5[222]; 
                dec[223] <= (a223_2 == 8'b0) & errs4 ? ~r5[223] : r5[223]; 
                dec[224] <= (a224_2 == 8'b0) & errs4 ? ~r5[224] : r5[224]; 
                dec[225] <= (a225_2 == 8'b0) & errs4 ? ~r5[225] : r5[225]; 
                dec[226] <= (a226_2 == 8'b0) & errs4 ? ~r5[226] : r5[226]; 
                dec[227] <= (a227_2 == 8'b0) & errs4 ? ~r5[227] : r5[227]; 
                dec[228] <= (a228_2 == 8'b0) & errs4 ? ~r5[228] : r5[228]; 
                dec[229] <= (a229_2 == 8'b0) & errs4 ? ~r5[229] : r5[229]; 
                dec[230] <= (a230_2 == 8'b0) & errs4 ? ~r5[230] : r5[230]; 
                dec[231] <= (a231_2 == 8'b0) & errs4 ? ~r5[231] : r5[231]; 
                dec[232] <= (a232_2 == 8'b0) & errs4 ? ~r5[232] : r5[232]; 
                dec[233] <= (a233_2 == 8'b0) & errs4 ? ~r5[233] : r5[233]; 
                dec[234] <= (a234_2 == 8'b0) & errs4 ? ~r5[234] : r5[234]; 
                dec[235] <= (a235_2 == 8'b0) & errs4 ? ~r5[235] : r5[235]; 
                dec[236] <= (a236_2 == 8'b0) & errs4 ? ~r5[236] : r5[236]; 
                dec[237] <= (a237_2 == 8'b0) & errs4 ? ~r5[237] : r5[237]; 
                dec[238] <= (a238_2 == 8'b0) & errs4 ? ~r5[238] : r5[238]; 
                dec[239] <= (a239_2 == 8'b0) & errs4 ? ~r5[239] : r5[239]; 
                dec[240] <= (a240_2 == 8'b0) & errs4 ? ~r5[240] : r5[240]; 
                dec[241] <= (a241_2 == 8'b0) & errs4 ? ~r5[241] : r5[241]; 
                dec[242] <= (a242_2 == 8'b0) & errs4 ? ~r5[242] : r5[242]; 
                dec[243] <= (a243_2 == 8'b0) & errs4 ? ~r5[243] : r5[243]; 
                dec[244] <= (a244_2 == 8'b0) & errs4 ? ~r5[244] : r5[244]; 
                dec[245] <= (a245_2 == 8'b0) & errs4 ? ~r5[245] : r5[245]; 
                dec[246] <= (a246_2 == 8'b0) & errs4 ? ~r5[246] : r5[246]; 
                dec[247] <= (a247_2 == 8'b0) & errs4 ? ~r5[247] : r5[247]; 
                dec[248] <= (a248_2 == 8'b0) & errs4 ? ~r5[248] : r5[248]; 
                dec[249] <= (a249_2 == 8'b0) & errs4 ? ~r5[249] : r5[249]; 
                dec[250] <= (a250_2 == 8'b0) & errs4 ? ~r5[250] : r5[250]; 
                dec[251] <= (a251_2 == 8'b0) & errs4 ? ~r5[251] : r5[251]; 
                dec[252] <= (a252_2 == 8'b0) & errs4 ? ~r5[252] : r5[252]; 
                dec[253] <= (a253_2 == 8'b0) & errs4 ? ~r5[253] : r5[253]; 
                dec[254] <= (a254_2 == 8'b0) & errs4 ? ~r5[254] : r5[254]; 
 


                dec[255] <= r5[255] ^ d_e;
//                dec[15] <= errs2 ? r3[15] ^ d_e : r3[15] ^ d_e ^ 1'b1;
            end else
                dec <= r5;
        
        end
    end
    
endmodule
