`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/02/2024 07:12:37 AM
// Design Name: 
// Module Name: PC_bsc_channel_block_ebch_256_239
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PC_bsc_channel_block_ebch_256_239(
    input clk,
    input reset,
    input wire [8191:0] seed,
    input wire [15:0] cross_prob,
    input  wire [255:0] codeword1,
    input  wire [255:0] codeword2,
    input  wire [255:0] codeword3,
    input  wire [255:0] codeword4,
    input  wire [255:0] codeword5,
    input  wire [255:0] codeword6,
    input  wire [255:0] codeword7,
    input  wire [255:0] codeword8,
    input  wire [255:0] codeword9,
    input  wire [255:0] codeword10,
    input  wire [255:0] codeword11,
    input  wire [255:0] codeword12,
    input  wire [255:0] codeword13,
    input  wire [255:0] codeword14,
    input  wire [255:0] codeword15,
    input  wire [255:0] codeword16,
    output wire  [255:0] received1,
    output wire  [255:0] received2,
    output wire  [255:0] received3,
    output wire  [255:0] received4,
    output wire  [255:0] received5,
    output wire  [255:0] received6,
    output wire  [255:0] received7,
    output wire  [255:0] received8,
    output wire  [255:0] received9,
    output wire  [255:0] received10,
    output wire  [255:0] received11,
    output wire  [255:0] received12,
    output wire  [255:0] received13,
    output wire  [255:0] received14,
    output wire  [255:0] received15,
    output wire  [255:0] received16
    );
    
//    reg [4095:0] seed1;
//    reg [4095:0] seed2;
//    reg [4095:0] seed3;
//    reg [4095:0] seed4;
//    reg [4095:0] seed5;
//    reg [4095:0] seed6;
//    reg [4095:0] seed7;
//    reg [4095:0] seed8;
//    reg [4095:0] seed9;
//    reg [4095:0] seed10;
//    reg [4095:0] seed11;
//    reg [4095:0] seed12;
//    reg [4095:0] seed13;
//    reg [4095:0] seed14;
//    reg [4095:0] seed15;
//    reg [4095:0] seed16;
    
//    always@ (posedge clk) begin
//        seed1 <= {seed[1227],seed[2508],seed[1106],seed[543],seed[3292],seed[2432],seed[1097],seed[2437],seed[1154],seed[1644],seed[3327],seed[1620],seed[25],seed[1404],seed[2426],seed[1993],seed[463],seed[2638],seed[2804],seed[671],seed[927],seed[3516],seed[54],seed[7],seed[859],seed[648],seed[2616],seed[2593],seed[2880],seed[3772],seed[1755],seed[2394],seed[2021],seed[2525],seed[2233],seed[2965],seed[2323],seed[3719],seed[2167],seed[143],seed[1652],seed[990],seed[1495],seed[1220],seed[75],seed[2570],seed[202],seed[2014],seed[3864],seed[3013],seed[3214],seed[1998],seed[2296],seed[532],seed[523],seed[379],seed[3116],seed[1668],seed[1746],seed[695],seed[490],seed[3887],seed[3315],seed[2571],seed[3671],seed[3740],seed[2254],seed[1735],seed[1113],seed[2645],seed[1301],seed[23],seed[460],seed[253],seed[186],seed[3471],seed[3979],seed[893],seed[3350],seed[3570],seed[2642],seed[4056],seed[1233],seed[2791],seed[3421],seed[913],seed[2294],seed[158],seed[3794],seed[2895],seed[3591],seed[3764],seed[779],seed[1364],seed[4026],seed[3910],seed[3991],seed[218],seed[541],seed[1198],seed[3127],seed[1088],seed[670],seed[3707],seed[4086],seed[1875],seed[1325],seed[144],seed[2757],seed[113],seed[4054],seed[3607],seed[1509],seed[3282],seed[2382],seed[1419],seed[2983],seed[2482],seed[185],seed[1247],seed[2255],seed[1833],seed[1855],seed[615],seed[1557],seed[896],seed[3766],seed[1276],seed[2594],seed[562],seed[1929],seed[3807],seed[3852],seed[2524],seed[3552],seed[832],seed[3551],seed[2654],seed[940],seed[678],seed[2991],seed[276],seed[1067],seed[833],seed[1210],seed[3657],seed[888],seed[2945],seed[427],seed[3658],seed[3654],seed[3232],seed[898],seed[3435],seed[3888],seed[593],seed[518],seed[433],seed[3799],seed[660],seed[2690],seed[3099],seed[2583],seed[3792],seed[135],seed[169],seed[3999],seed[1902],seed[3021],seed[472],seed[1409],seed[3870],seed[1654],seed[3428],seed[181],seed[2313],seed[1188],seed[3086],seed[3128],seed[3094],seed[596],seed[232],seed[209],seed[3803],seed[3755],seed[2155],seed[3411],seed[2126],seed[1085],seed[2700],seed[2089],seed[2454],seed[340],seed[2213],seed[105],seed[3412],seed[2780],seed[96],seed[3083],seed[3381],seed[3631],seed[2451],seed[3301],seed[1141],seed[4042],seed[2103],seed[1104],seed[2678],seed[1546],seed[3082],seed[2116],seed[1624],seed[2694],seed[193],seed[2952],seed[3668],seed[2993],seed[2316],seed[3929],seed[2272],seed[821],seed[3268],seed[2201],seed[243],seed[1318],seed[1844],seed[617],seed[774],seed[819],seed[234],seed[2440],seed[439],seed[581],seed[527],seed[142],seed[1846],seed[2994],seed[1782],seed[134],seed[3366],seed[3946],seed[633],seed[2695],seed[1817],seed[569],seed[2207],seed[3394],seed[1921],seed[3944],seed[2276],seed[3811],seed[414],seed[509],seed[1870],seed[1759],seed[891],seed[422],seed[3859],seed[4],seed[466],seed[22],seed[822],seed[338],seed[3647],seed[3741],seed[2541],seed[2093],seed[1692],seed[2953],seed[3300],seed[2239],seed[1084],seed[1629],seed[2020],seed[1768],seed[2234],seed[3066],seed[2324],seed[281],seed[547],seed[634],seed[1825],seed[1293],seed[259],seed[520],seed[907],seed[1648],seed[97],seed[592],seed[2340],seed[1513],seed[174],seed[3734],seed[599],seed[2134],seed[2724],seed[1878],seed[2259],seed[3016],seed[3360],seed[1882],seed[291],seed[761],seed[428],seed[199],seed[628],seed[1715],seed[872],seed[1248],seed[2794],seed[407],seed[843],seed[2297],seed[3841],seed[3050],seed[279],seed[2310],seed[2264],seed[1723],seed[3184],seed[2876],seed[957],seed[3011],seed[842],seed[1436],seed[1559],seed[3438],seed[91],seed[2899],seed[2359],seed[180],seed[3558],seed[692],seed[258],seed[1476],seed[3917],seed[533],seed[2919],seed[3409],seed[1699],seed[1549],seed[1359],seed[1566],seed[2623],seed[3873],seed[3364],seed[2399],seed[1612],seed[3642],seed[3244],seed[392],seed[1901],seed[3967],seed[2818],seed[2946],seed[2352],seed[4091],seed[1679],seed[99],seed[1693],seed[1724],seed[2085],seed[1795],seed[398],seed[13],seed[231],seed[70],seed[3565],seed[1616],seed[2712],seed[487],seed[1398],seed[1353],seed[580],seed[4043],seed[1203],seed[489],seed[94],seed[840],seed[1176],seed[2607],seed[1029],seed[3156],seed[2873],seed[3203],seed[3983],seed[2446],seed[1414],seed[3957],seed[3447],seed[2867],seed[2223],seed[3492],seed[221],seed[1574],seed[2447],seed[3208],seed[3371],seed[29],seed[924],seed[3238],seed[133],seed[3161],seed[3387],seed[3950],seed[673],seed[1063],seed[3400],seed[2337],seed[3532],seed[697],seed[4068],seed[519],seed[1142],seed[1390],seed[1206],seed[1927],seed[3786],seed[4012],seed[557],seed[3334],seed[2245],seed[1886],seed[3056],seed[2069],seed[3134],seed[2145],seed[2746],seed[735],seed[2051],seed[2733],seed[81],seed[3789],seed[2332],seed[2626],seed[3470],seed[192],seed[227],seed[1773],seed[368],seed[1776],seed[1584],seed[920],seed[2606],seed[720],seed[3678],seed[1893],seed[3049],seed[1861],seed[1308],seed[2148],seed[828],seed[2967],seed[3320],seed[3069],seed[1483],seed[1672],seed[3927],seed[2424],seed[84],seed[3940],seed[3380],seed[1591],seed[2956],seed[892],seed[1857],seed[1610],seed[665],seed[1134],seed[986],seed[3439],seed[528],seed[1568],seed[2665],seed[3397],seed[900],seed[1479],seed[1722],seed[1767],seed[330],seed[1634],seed[1055],seed[3129],seed[3098],seed[1137],seed[1852],seed[1830],seed[2331],seed[3197],seed[3425],seed[2811],seed[3237],seed[3540],seed[383],seed[2191],seed[1018],seed[1793],seed[2681],seed[118],seed[3589],seed[3302],seed[1373],seed[2787],seed[2820],seed[4009],seed[2256],seed[352],seed[2403],seed[3923],seed[213],seed[559],seed[654],seed[1529],seed[3499],seed[4011],seed[1347],seed[4030],seed[3667],seed[2640],seed[984],seed[864],seed[579],seed[1717],seed[1528],seed[2909],seed[1785],seed[2949],seed[1482],seed[1384],seed[2793],seed[1408],seed[2664],seed[1897],seed[3026],seed[3939],seed[1499],seed[3139],seed[1473],seed[2462],seed[709],seed[1057],seed[611],seed[813],seed[1514],seed[3234],seed[3406],seed[2326],seed[1845],seed[1681],seed[2035],seed[2227],seed[3462],seed[384],seed[1890],seed[2445],seed[434],seed[3229],seed[2158],seed[825],seed[2796],seed[2822],seed[1311],seed[582],seed[1895],seed[1771],seed[3006],seed[2527],seed[139],seed[3575],seed[3079],seed[928],seed[2932],seed[851],seed[1952],seed[3716],seed[1205],seed[146],seed[385],seed[3791],seed[2143],seed[2305],seed[155],seed[469],seed[4064],seed[3919],seed[3801],seed[59],seed[788],seed[3963],seed[1928],seed[537],seed[3655],seed[542],seed[722],seed[3324],seed[2773],seed[2137],seed[3812],seed[223],seed[2784],seed[3624],seed[1996],seed[1385],seed[3926],seed[3760],seed[576],seed[1918],seed[2749],seed[393],seed[2769],seed[1268],seed[2772],seed[3019],seed[3553],seed[3456],seed[3988],seed[2529],seed[734],seed[2622],seed[1179],seed[3797],seed[2418],seed[175],seed[4093],seed[979],seed[1617],seed[1659],seed[1696],seed[3603],seed[1209],seed[3871],seed[1963],seed[2173],seed[2037],seed[1147],seed[2885],seed[103],seed[626],seed[3109],seed[3287],seed[2697],seed[2986],seed[3351],seed[1037],seed[2419],seed[436],seed[1231],seed[2829],seed[3155],seed[555],seed[3533],seed[2483],seed[1302],seed[3866],seed[1753],seed[1274],seed[1791],seed[621],seed[195],seed[587],seed[172],seed[3115],seed[1031],seed[3095],seed[3259],seed[170],seed[1720],seed[961],seed[1335],seed[1238],seed[1687],seed[1118],seed[3555],seed[3040],seed[2217],seed[3643],seed[4065],seed[3133],seed[1333],seed[3976],seed[1994],seed[306],seed[3293],seed[1326],seed[2547],seed[1619],seed[2591],seed[4057],seed[3121],seed[403],seed[3105],seed[3077],seed[72],seed[3557],seed[2628],seed[1809],seed[1168],seed[2834],seed[1937],seed[3452],seed[298],seed[2280],seed[2864],seed[3977],seed[3507],seed[2457],seed[1639],seed[246],seed[1818],seed[2602],seed[3503],seed[2067],seed[3743],seed[343],seed[1805],seed[2955],seed[2709],seed[753],seed[1425],seed[2146],seed[4017],seed[3189],seed[3487],seed[2325],seed[2110],seed[1540],seed[77],seed[3955],seed[1623],seed[3501],seed[3691],seed[2329],seed[3297],seed[3612],seed[2542],seed[4031],seed[1224],seed[3329],seed[3619],seed[566],seed[981],seed[1292],seed[121],seed[855],seed[2463],seed[4069],seed[3855],seed[2514],seed[2611],seed[3442],seed[723],seed[3798],seed[3395],seed[409],seed[1050],seed[2963],seed[1920],seed[2226],seed[3266],seed[1820],seed[2376],seed[3878],seed[1675],seed[1530],seed[2655],seed[442],seed[3032],seed[3247],seed[1502],seed[2502],seed[1150],seed[2300],seed[431],seed[3845],seed[3554],seed[1126],seed[3393],seed[1757],seed[2420],seed[2790],seed[1339],seed[3308],seed[705],seed[2806],seed[4052],seed[3168],seed[870],seed[3340],seed[1489],seed[1831],seed[4010],seed[3010],seed[3354],seed[2472],seed[1816],seed[3769],seed[2471],seed[1064],seed[110],seed[2357],seed[1909],seed[3055],seed[326],seed[3463],seed[295],seed[2507],seed[1307],seed[2936],seed[2042],seed[3973],seed[1058],seed[3166],seed[2598],seed[1714],seed[3593],seed[1321],seed[288],seed[2910],seed[539],seed[1520],seed[2208],seed[2004],seed[755],seed[1880],seed[680],seed[737],seed[3971],seed[3728],seed[2595],seed[2624],seed[2795],seed[3294],seed[3722],seed[1131],seed[553],seed[1285],seed[1907],seed[3724],seed[1941],seed[3897],seed[63],seed[3446],seed[701],seed[3997],seed[1556],seed[1636],seed[2985],seed[922],seed[650],seed[3260],seed[2676],seed[1152],seed[359],seed[2517],seed[1740],seed[353],seed[3020],seed[1627],seed[1704],seed[2520],seed[3907],seed[1649],seed[827],seed[1],seed[1609],seed[2609],seed[2816],seed[560],seed[3171],seed[2923],seed[1066],seed[1146],seed[911],seed[2815],seed[2738],seed[222],seed[1484],seed[1194],seed[3090],seed[2835],seed[2405],seed[1637],seed[770],seed[18],seed[1498],seed[1277],seed[767],seed[2311],seed[2767],seed[3683],seed[959],seed[205],seed[1362],seed[1047],seed[1828],seed[3521],seed[2629],seed[2212],seed[4040],seed[2088],seed[488],seed[885],seed[880],seed[980],seed[1580],seed[1647],seed[3935],seed[2590],seed[3508],seed[4087],seed[21],seed[3602],seed[196],seed[3932],seed[1433],seed[263],seed[563],seed[1177],seed[71],seed[3306],seed[1181],seed[3833],seed[3617],seed[2358],seed[1738],seed[3851],seed[292],seed[3921],seed[2289],seed[3249],seed[3213],seed[3087],seed[2801],seed[3182],seed[948],seed[405],seed[2027],seed[458],seed[1618],seed[1402],seed[4001],seed[610],seed[173],seed[1242],seed[1173],seed[3776],seed[1374],seed[2417],seed[1167],seed[3609],seed[3633],seed[3410],seed[974],seed[1917],seed[43],seed[2371],seed[1239],seed[2006],seed[3399],seed[2854],seed[3365],seed[3111],seed[2287],seed[381],seed[1216],seed[1544],seed[2355],seed[1581],seed[651],seed[3423],seed[416],seed[2937],seed[201],seed[93],seed[1615],seed[2969],seed[884],seed[3699],seed[1972],seed[2778],seed[2905],seed[3547],seed[2637],seed[2900],seed[2029],seed[3067],seed[3818],seed[3781],seed[2238],seed[3538],seed[661],seed[903],seed[3120],seed[797],seed[2510],seed[516],seed[3649],seed[360],seed[3909],seed[2001],seed[2277],seed[2040],seed[2762],seed[37],seed[3536],seed[1430],seed[3641],seed[1606],seed[1105],seed[2842],seed[1368],seed[4049],seed[2914],seed[1829],seed[423],seed[334],seed[117],seed[3383],seed[2858],seed[305],seed[4021],seed[3341],seed[3960],seed[841],seed[848],seed[3088],seed[1564],seed[679],seed[3338],seed[1860],seed[3986],seed[1748],seed[2187],seed[2667],seed[852],seed[3714],seed[507],seed[2597],seed[983],seed[3860],seed[3648],seed[130],seed[991],seed[2281],seed[1132],seed[2002],seed[255],seed[534],seed[20],seed[415],seed[3241],seed[1367],seed[1572],seed[718],seed[2828],seed[1447],seed[1360],seed[623],seed[3632],seed[3479],seed[787],seed[2916],seed[1645],seed[2630],seed[402],seed[2050],seed[1014],seed[785],seed[244],seed[2041],seed[2232],seed[2209],seed[491],seed[600],seed[782],seed[3936],seed[877],seed[760],seed[3461],seed[830],seed[3636],seed[1613],seed[1267],seed[1261],seed[2430],seed[696],seed[24],seed[260],seed[3690],seed[2499],seed[784],seed[2074],seed[741],seed[3024],seed[2468],seed[2601],seed[1330],seed[607],seed[3257],seed[3543],seed[283],seed[3753],seed[2887],seed[824],seed[1832],seed[2269],seed[2282],seed[2071],seed[3968],seed[742],seed[3071],seed[2157],seed[4006],seed[3969],seed[2713],seed[3408],seed[3686],seed[3842],seed[3065],seed[2328],seed[3829],seed[2200],seed[1211],seed[1357],seed[3018],seed[2861],seed[3003],seed[1734],seed[875],seed[3858],seed[1464],seed[1036],seed[1600],seed[2079],seed[40],seed[357],seed[3726],seed[4051],seed[3415],seed[1640],seed[3583],seed[4039],seed[1604],seed[814],seed[86],seed[3359],seed[854],seed[2843],seed[2911],seed[2260],seed[895],seed[2068],seed[1543],seed[2125],seed[2917],seed[2719],seed[646],seed[3270],seed[411],seed[1913],seed[938],seed[3494],seed[1579],seed[3809],seed[1096],seed[1287],seed[2752],seed[1388],seed[776],seed[1685],seed[3820],seed[1349],seed[1243],seed[2696],seed[2689],seed[1822],seed[2947],seed[3110],seed[881],seed[3418],seed[1214],seed[2186],seed[2774],seed[2679],seed[120],seed[2935],seed[3186],seed[2295],seed[1991],seed[3837],seed[2604],seed[1281],seed[2896],seed[1578],seed[733],seed[1790],seed[597],seed[3332],seed[1924],seed[1166],seed[4008],seed[3763],seed[1719],seed[1800],seed[2485],seed[2763],seed[2028],seed[1823],seed[479],seed[311],seed[603],seed[2240],seed[1508],seed[1827],seed[1742],seed[2782],seed[2384],seed[2727],seed[750],seed[3272],seed[1475],seed[3075],seed[1710],seed[3510],seed[441],seed[3876],seed[2686],seed[2308],seed[548],seed[1417],seed[2580],seed[769],seed[2532],seed[1535],seed[2109],seed[883],seed[3254],seed[1487],seed[2924],seed[128],seed[3243],seed[1560],seed[3444],seed[3250],seed[1836],seed[3277],seed[2195],seed[1080],seed[530],seed[1872],seed[3738],seed[627],seed[3634],seed[1076],seed[4025],seed[3422],seed[325],seed[1966],seed[3312],seed[1807],seed[2474],seed[1550],seed[3942],seed[1413],seed[2488],seed[745],seed[2996],seed[3046],seed[3718],seed[823],seed[585],seed[1752],seed[2734],seed[2184],seed[996],seed[1102],seed[4090],seed[2587],seed[3022],seed[3504],seed[2284],seed[2242],seed[1159],seed[3937],seed[987],seed[2862],seed[3733],seed[200],seed[3568],seed[1418],seed[3822],seed[1571],seed[1423],seed[3262],seed[480],seed[1949],seed[1303],seed[951],seed[282],seed[2064],seed[638],seed[2120],seed[2177],seed[4078],seed[1984],seed[316],seed[1358],seed[1389],seed[3037],seed[1381],seed[2721],seed[2731],seed[3154],seed[2224],seed[3588],seed[2891],seed[3629],seed[2452],seed[1300],seed[2768],seed[125],seed[64],seed[275],seed[3879],seed[3677],seed[3981],seed[3458],seed[3891],seed[1200],seed[2631],seed[3443],seed[52],seed[937],seed[304],seed[1053],seed[3496],seed[740],seed[2617],seed[2559],seed[80],seed[1938],seed[3062],seed[2270],seed[3373],seed[3747],seed[1153],seed[1183],seed[1437],seed[484],seed[588],seed[485],seed[4083],seed[2106],seed[2258],seed[2022],seed[1270],seed[656],seed[450],seed[1298],seed[529],seed[946],seed[167],seed[2391],seed[3271],seed[2298],seed[3356],seed[1077],seed[157],seed[2564],seed[2176],seed[3303],seed[2663],seed[1932],seed[3759],seed[3137],seed[0],seed[4070],seed[3],seed[449],seed[1427],seed[1667],seed[3468],seed[693],seed[2135],seed[2342],seed[207],seed[2413],seed[438],seed[1288],seed[3836],seed[2644],seed[1943],seed[3651],seed[2132],seed[1934],seed[2929],seed[274],seed[1232],seed[2379],seed[371],seed[1324],seed[1174],seed[2897],seed[1967],seed[2855],seed[1987],seed[3500],seed[3033],seed[1497],seed[3795],seed[2660],seed[1485],seed[2839],seed[2012],seed[3188],seed[3542],seed[2797],seed[2693],seed[3138],seed[3124],seed[2530],seed[2668],seed[1968],seed[1631],seed[932],seed[3093],seed[1969],seed[1350],seed[3278],seed[2998],seed[3349],seed[49],seed[214],seed[1850],seed[287],seed[1910],seed[3353],seed[1980],seed[2222],seed[2097],seed[210],seed[313],seed[2692],seed[224],seed[254],seed[3779],seed[1607],seed[3289],seed[3611],seed[3190],seed[2343],seed[3523],seed[690],seed[3970],seed[3497],seed[3073],seed[1130],seed[1702],seed[3592],seed[3493],seed[1611],seed[2557],seed[1678],seed[567],seed[2531],seed[2312],seed[290],seed[794],seed[982],seed[1810],seed[335],seed[1554],seed[2671],seed[796],seed[448],seed[1576],seed[2129],seed[3343],seed[2632],seed[2776],seed[577],seed[905],seed[3846],seed[4033],seed[2206],seed[3625],seed[3665],seed[150],seed[2330],seed[2438],seed[3585],seed[2095],seed[775],seed[3346],seed[3265],seed[406],seed[3347],seed[2718],seed[3159],seed[236],seed[916],seed[879],seed[3160],seed[1835],seed[1240],seed[1582],seed[1124],seed[3377],seed[2893],seed[2180],seed[219],seed[3001],seed[2183],seed[1575],seed[376],seed[2560],seed[1628],seed[3034],seed[1555],seed[2511],seed[1745],seed[1143],seed[3739],seed[417],seed[2056],seed[332],seed[3512],seed[554],seed[3045],seed[2883],seed[272],seed[2526],seed[4082],seed[358],seed[41],seed[3404],seed[2464],seed[2741],seed[4036],seed[2698],seed[453],seed[3749],seed[2049],seed[1761],seed[2759],seed[2901],seed[3267],seed[2725],seed[3630],seed[2387],seed[2026],seed[3194],seed[754],seed[2652],seed[2860],seed[3054],seed[1445],seed[3574],seed[3783],seed[1098],seed[267],seed[2516],seed[2119],seed[2484],seed[2107],seed[1521],seed[38],seed[866],seed[1492],seed[3269],seed[1320],seed[871],seed[389],seed[3273],seed[849],seed[2404],seed[2980],seed[296],seed[1565],seed[129],seed[2573],seed[16],seed[1283],seed[2635],seed[3118],seed[3616],seed[772],seed[2214],seed[853],seed[2024],seed[2651],seed[3736],seed[799],seed[3948],seed[2203],seed[2549],seed[319],seed[918],seed[252],seed[1586],seed[3370],seed[1252],seed[399],seed[437],seed[418],seed[1762],seed[2388],seed[771],seed[257],seed[2202],seed[3587],seed[1990],seed[1597],seed[2925],seed[1208],seed[3610],seed[3474],seed[1510],seed[3117],seed[978],seed[2467],seed[1642],seed[1093],seed[1501],seed[2052],seed[2448],seed[1455],seed[2096],seed[2370],seed[3869],seed[467],seed[3793],seed[3990],seed[2934],seed[1415],seed[2309],seed[3951],seed[3417],seed[3582],seed[882],seed[2592],seed[2179],seed[2962],seed[2237],seed[3815],seed[2892],seed[1522],seed[4095],seed[1770],seed[92],seed[1079],seed[455],seed[1854],seed[1100],seed[684],seed[2603],seed[1989],seed[2981],seed[2904],seed[2303],seed[934],seed[1392],seed[2301],seed[3255],seed[570],seed[1016],seed[1518],seed[1013],seed[1361],seed[2657],seed[3908],seed[1295],seed[2423],seed[2154],seed[1786],seed[1022],seed[2299],seed[668],seed[3701],seed[3856],seed[2216],seed[3051],seed[2168],seed[1342],seed[2252],seed[886],seed[3389],seed[1226],seed[1673],seed[3429],seed[909],seed[565],seed[2378],seed[944],seed[2572],seed[1467],seed[2821],seed[2008],seed[1784],seed[347],seed[369],seed[3502],seed[208],seed[3078],seed[1657],seed[1733],seed[2722],seed[61],seed[746],seed[2827],seed[1806],seed[837],seed[3113],seed[1906],seed[942],seed[874],seed[688],seed[2519],seed[1397],seed[1383],seed[3176],seed[3644],seed[3092],seed[3455],seed[2112],seed[2372],seed[1365],seed[2605],seed[3295],seed[2480],seed[3674],seed[1470],seed[2555],seed[85],seed[2044],seed[1936],seed[575],seed[3276],seed[459],seed[3027],seed[2427],seed[1382],seed[2845],seed[156],seed[598],seed[2927],seed[1466],seed[3253],seed[3645],seed[1780],seed[1663],seed[2215],seed[12],seed[618],seed[3918],seed[2118],seed[3322],seed[171],seed[1834],seed[3169],seed[56],seed[3445],seed[127],seed[3883],seed[2491],seed[2374],seed[1289],seed[2755],seed[8],seed[477],seed[413],seed[395],seed[624],seed[3985],seed[1265],seed[925],seed[154],seed[2055],seed[1869],seed[3828],seed[3331],seed[1935],seed[2979],seed[1481],seed[1655],seed[3806],seed[1751],seed[2381],seed[2278],seed[3219],seed[3752],seed[35],seed[3486],seed[613],seed[1337],seed[2128],seed[2354],seed[1109],seed[44],seed[1876],seed[998],seed[3344],seed[672],seed[4028],seed[2817],seed[2481],seed[1279],seed[1838],seed[27],seed[3785],seed[3835],seed[730],seed[1690],seed[309],seed[229],seed[2569],seed[2494],seed[1428],seed[3060],seed[3770],seed[230],seed[3639],seed[1898],seed[635],seed[114],seed[1212],seed[1336],seed[3978],seed[1983],seed[1169],seed[2477],seed[2150],seed[3672],seed[2080],seed[1553],seed[3717],seed[3142],seed[2961],seed[1879],seed[1658],seed[1865],seed[1905],seed[1450],seed[166],seed[2879],seed[710],seed[1567],seed[1583],seed[107],seed[1904],seed[1848],seed[2000],seed[2091],seed[3653],seed[2496],seed[2868],seed[2218],seed[2105],seed[1222],seed[1551],seed[2959],seed[3070],seed[969],seed[2551],seed[65],seed[3059],seed[106],seed[4059],seed[3945],seed[2992],seed[1074],seed[1766],seed[3413],seed[159],seed[2761],seed[1376],seed[2705],seed[3546],seed[2523],seed[1352],seed[2025],seed[1587],seed[4060],seed[57],seed[447],seed[34],seed[3029],seed[1725],seed[2383],seed[1033],seed[2841],seed[3482],seed[492],seed[3802],seed[2136],seed[3920],seed[3367],seed[2365],seed[3164],seed[3566],seed[3576],seed[2409],seed[2063],seed[1228],seed[2054],seed[67],seed[2625],seed[873],seed[3431],seed[2100],seed[3434],seed[3426],seed[3089],seed[867],seed[1071],seed[708],seed[985],seed[493],seed[2972],seed[504],seed[198],seed[1396],seed[3775],seed[2938],seed[1900],seed[1930],seed[2034],seed[3158],seed[3721],seed[876],seed[939],seed[564],seed[2647],seed[4007],seed[3746],seed[1032],seed[4089],seed[1442],seed[3601],seed[3025],seed[1314],seed[1923],seed[2402],seed[3572],seed[3831],seed[977],seed[3200],seed[2416],seed[1117],seed[1743],seed[2706],seed[540],seed[4050],seed[2369],seed[3378],seed[3626],seed[112],seed[1813],seed[1044],seed[248],seed[2567],seed[2509],seed[1674],seed[686],seed[691],seed[1970],seed[2292],seed[2009],seed[400],seed[496],seed[2826],seed[3005],seed[1925],seed[1887],seed[3898],seed[1729],seed[1812],seed[2246],seed[445],seed[2673],seed[2196],seed[1940],seed[950],seed[3074],seed[715],seed[4032],seed[2585],seed[1123],seed[3449],seed[2401],seed[2926],seed[857],seed[4023],seed[2730],seed[2831],seed[1056],seed[3141],seed[3012],seed[1371],seed[2521],seed[1908],seed[1682],seed[3192],seed[816],seed[3635],seed[2077],seed[2715],seed[926],seed[4081],seed[666],seed[2639],seed[2613],seed[3790],seed[3205],seed[747],seed[310],seed[1230],seed[4080],seed[3638],seed[2850],seed[674],seed[820],seed[1533],seed[1051],seed[3628],seed[4074],seed[1468],seed[153],seed[1421],seed[3526],seed[2265],seed[639],seed[3682],seed[1331],seed[1394],seed[1027],seed[2273],seed[2141],seed[62],seed[3152],seed[2373],seed[887],seed[2266],seed[869],seed[3949],seed[2497],seed[2030],seed[151],seed[2503],seed[2680],seed[126],seed[3467],seed[3044],seed[1236],seed[2500],seed[277],seed[131],seed[1244],seed[3476],seed[1792],seed[2353],seed[3505],seed[1922],seed[240],seed[1781],seed[2957],seed[268],seed[1511],seed[994],seed[2288],seed[2364],seed[3750],seed[2243],seed[2770],seed[2348],seed[2728],seed[804],seed[3123],seed[1278],seed[1662],seed[2389],seed[1945],seed[764],seed[3398],seed[3915],seed[3998],seed[815],seed[375],seed[3995],seed[1758],seed[3847],seed[3352],seed[1234],seed[3202],seed[464],seed[1112],seed[963],seed[2977],seed[1387],seed[3854],seed[3085],seed[1840],seed[3256],seed[3788],seed[2247],seed[2674],seed[2],seed[3311],seed[1976],seed[1665],seed[1814],seed[3709],seed[2575],seed[3135],seed[3737],seed[2964],seed[1115],seed[3615],seed[474],seed[2669],seed[2410],seed[3913],seed[675],seed[109],seed[1457],seed[526],seed[2837],seed[1175],seed[2533],seed[1089],seed[2720],seed[391],seed[3107],seed[1633],seed[2600],seed[846],seed[3531],seed[2553],seed[780],seed[2013],seed[3901],seed[3596],seed[2094],seed[1237],seed[2918],seed[2648],seed[3436],seed[3982],seed[2479],seed[719],seed[3966],seed[1120],seed[2807],seed[3843],seed[2138],seed[3172],seed[2833],seed[204],seed[2458],seed[1161],seed[410],seed[1561],seed[2274],seed[152],seed[2019],seed[1709],seed[3405],seed[3796],seed[3535],seed[707],seed[1266],seed[4075],seed[988],seed[1221],seed[1802],seed[1730],seed[972],seed[115],seed[1635],seed[2475],seed[2701],seed[2211],seed[1862],seed[1400],seed[3757],seed[952],seed[3206],seed[3685],seed[2059],seed[2115],seed[3207],seed[2775],seed[2251],seed[68],seed[2554],seed[3577],seed[315],seed[2812],seed[2033],seed[751],seed[1165],seed[3209],seed[2408],seed[706],seed[362],seed[2320],seed[233],seed[2263],seed[3545],seed[3830],seed[1946],seed[1107],seed[2318],seed[265],seed[2459],seed[2687],seed[3102],seed[3170],seed[2181],seed[2267],seed[2130],seed[1892],seed[2236],seed[714],seed[1703],seed[1839],seed[1046],seed[2546],seed[2261],seed[3893],seed[1092],seed[271],seed[968],seed[3882],seed[30],seed[187],seed[1191],seed[954],seed[1598],seed[1005],seed[1939],seed[1386],seed[2851],seed[1988],seed[3047],seed[4037],seed[3827],seed[264],seed[1125],seed[4055],seed[1081],seed[3149],seed[971],seed[235],seed[1821],seed[3711],seed[3742],seed[184],seed[1552],seed[1128],seed[3491],seed[1926],seed[478],seed[2073],seed[1114],seed[2166],seed[2087],seed[3038],seed[2920],seed[2053],seed[4016],seed[3961],seed[1355],seed[643],seed[2522],seed[162],seed[1344],seed[1465],seed[2174],seed[2058],seed[2810],seed[862],seed[1916],seed[73],seed[3787],seed[3941],seed[11],seed[3911],seed[2043],seed[1585],seed[2888],seed[1819],seed[1171],seed[2726],seed[2439],seed[1315],seed[3895],seed[732],seed[495],seed[1997],seed[468],seed[752],seed[2171],seed[1708],seed[834],seed[331],seed[1217],seed[1646],seed[237],seed[1894],seed[1195],seed[462],seed[440],seed[2205],seed[552],seed[676],seed[3586],seed[793],seed[404],seed[2066],seed[3178],seed[3224],seed[960],seed[1170],seed[486],seed[2487],seed[3824],seed[1779],seed[3490],seed[2661],seed[2133],seed[1193],seed[1023],seed[2544],seed[2341],seed[1182],seed[658],seed[1537],seed[2881],seed[501],seed[66],seed[2513],seed[572],seed[1853],seed[3825],seed[653],seed[344],seed[3333],seed[3361],seed[3745],seed[2460],seed[3126],seed[3725],seed[1269],seed[3488],seed[1688],seed[1446],seed[2743],seed[749],seed[931],seed[3153],seed[2380],seed[1933],seed[3305],seed[102],seed[1348],seed[2235],seed[3771],seed[3280],seed[685],seed[1004],seed[2345],seed[1877],seed[1593],seed[3345],seed[3286],seed[1866],seed[1769],seed[1680],seed[763],seed[583],seed[3618],seed[420],seed[2366],seed[2204],seed[1523],seed[1881],seed[818],seed[3661],seed[3225],seed[2377],seed[2562],seed[289],seed[901],seed[2436],seed[3459],seed[3692],seed[3336],seed[1496],seed[1975],seed[179],seed[3712],seed[1366],seed[1911],seed[3518],seed[910],seed[3903],seed[2675],seed[1178],seed[3506],seed[1884],seed[682],seed[861],seed[3804],seed[3106],seed[1042],seed[728],seed[3465],seed[1562],seed[783],seed[2906],seed[1889],seed[836],seed[1686],seed[1858],seed[2540],seed[2392],seed[168],seed[293],seed[3819],seed[124],seed[3198],seed[1622],seed[844],seed[2007],seed[574],seed[620],seed[312],seed[2866],seed[3868],seed[811],seed[285],seed[372],seed[2225],seed[2882],seed[2819],seed[206],seed[1160],seed[2321],seed[3328],seed[1189],seed[2688],seed[2160],seed[941],seed[1985],seed[713],seed[1316],seed[3778],seed[808],seed[947],seed[3663],seed[147],seed[299],seed[2646],seed[1641],seed[294],seed[3478],seed[1590],seed[3342],seed[3623],seed[2621],seed[203],seed[3177],seed[88],seed[3689],seed[1973],seed[2199],seed[83],seed[4048],seed[3666],seed[3974],seed[3758],seed[2147],seed[777],seed[2090],seed[87],seed[1999],seed[663],seed[1246],seed[3727],seed[1062],seed[3520],seed[1713],seed[546],seed[374],seed[2633],seed[95],seed[1258],seed[894],seed[531],seed[3240],seed[2933],seed[1558],seed[100],seed[738],seed[3890],seed[602],seed[1180],seed[863],seed[970],seed[995],seed[1328],seed[2849],seed[2518],seed[1532],seed[3777],seed[1393],seed[2886],seed[2931],seed[2528],seed[3605],seed[3464],seed[3368],seed[3865],seed[538],seed[2512],seed[242],seed[3627],seed[1977],seed[3599],seed[2968],seed[161],seed[2290],seed[3580],seed[3216],seed[2971],seed[3402],seed[2162],seed[339],seed[1327],seed[3009],seed[1006],seed[3433],seed[3480],seed[1515],seed[4035],seed[2250],seed[3119],seed[2036],seed[1135],seed[2262],seed[2997],seed[2871],seed[1506],seed[3684],seed[182],seed[1061],seed[1797],seed[1486],seed[1136],seed[1015],seed[3659],seed[1341],seed[2574],seed[917],seed[2017],seed[9],seed[3251],seed[2170],seed[2057],seed[2443],seed[976],seed[2065],seed[1354],seed[1488],seed[3881],seed[845],seed[2039],seed[4015],seed[1859],seed[3773],seed[2102],seed[790],seed[524],seed[1025],seed[3076],seed[657],seed[3573],seed[997],seed[662],seed[1249],seed[3372],seed[435],seed[3097],seed[4047],seed[3556],seed[3309],seed[3813],seed[3694],seed[498],seed[3475],seed[3703],seed[1070],seed[1461],seed[1313],seed[1747],seed[1363],seed[3756],seed[386],seed[1961],seed[2407],seed[55],seed[2543],seed[739],seed[2393],seed[3840],seed[3637],seed[3564],seed[3730],seed[3140],seed[457],seed[256],seed[878],seed[625],seed[1028],seed[426],seed[2390],seed[999],seed[1286],seed[4071],seed[266],seed[3762],seed[3386],seed[380],seed[2535],seed[4077],seed[2178],seed[1040],seed[1202],seed[2588],seed[3191],seed[3581],seed[432],seed[545],seed[3318],seed[1503],seed[42],seed[1538],seed[2942],seed[1111],seed[2275],seed[1841],seed[2536],seed[3039],seed[2349],seed[101],seed[1103],seed[2940],seed[1660],seed[1312],seed[3004],seed[1605],seed[1694],seed[2060],seed[1959],seed[3290],seed[3590],seed[4002],seed[378],seed[317],seed[1643],seed[1405],seed[3880],seed[1356],seed[2156],seed[792],seed[3385],seed[2414],seed[1737],seed[3875],seed[3245],seed[3002],seed[614],seed[1669],seed[2185],seed[664],seed[558],seed[2677],seed[2431],seed[2608],seed[3849],seed[388],seed[1219],seed[2197],seed[3906],seed[3650],seed[2771],seed[2872],seed[3008],seed[3220],seed[762],seed[2825],seed[2003],seed[1676],seed[966],seed[2283],seed[1653],seed[3992],seed[341],seed[1625],seed[3481],seed[3183],seed[1749],seed[1218],seed[2104],seed[2747],seed[226],seed[4022],seed[1151],seed[1420],seed[2515],seed[3548],seed[3130],seed[3472],seed[4067],seed[3028],seed[3157],seed[2465],seed[51],seed[2078],seed[3620],seed[1310],seed[262],seed[1213],seed[2489],seed[2221],seed[2534],seed[3239],seed[3041],seed[3702],seed[1948],seed[342],seed[3061],seed[3030],seed[2010],seed[2788],seed[3321],seed[1411],seed[2350],seed[3103],seed[2783],seed[1078],seed[3457],seed[145],seed[3621],seed[616],seed[3180],seed[801],seed[2941],seed[1500],seed[3867],seed[3357],seed[3930],seed[1888],seed[322],seed[3477],seed[1319],seed[3195],seed[3081],seed[1626],seed[2113],seed[1808],seed[3780],seed[515],seed[3989],seed[647],seed[2466],seed[1458],seed[681],seed[3544],seed[550],seed[1577],seed[1589],seed[3165],seed[640],seed[2492],seed[2307],seed[4094],seed[953],seed[2684],seed[3122],seed[2636],seed[2153],seed[1187],seed[301],seed[1144],seed[2982],seed[1451],seed[3765],seed[2578],seed[1986],seed[2375],seed[280],seed[1121],seed[3975],seed[1273],seed[3104],seed[3928],seed[1684],seed[1380],seed[1811],seed[3705],seed[3330],seed[2428],seed[2581],seed[286],seed[1329],seed[2476],seed[3136],seed[2903],seed[3511],seed[3227],seed[703],seed[506],seed[1020],seed[2970],seed[250],seed[3774],seed[2351],seed[4005],seed[3108],seed[3660],seed[1095],seed[3844],seed[908],seed[2915],seed[2188],seed[2398],seed[2599],seed[1596],seed[328],seed[2169],seed[183],seed[3515],seed[3838],seed[1525],seed[2803],seed[2857],seed[4024],seed[3187],seed[3035],seed[1343],seed[4034],seed[212],seed[1410],seed[1296],seed[3112],seed[2335],seed[1192],seed[3369],seed[3744],seed[2415],seed[1241],seed[2228],seed[3222],seed[3114],seed[689],seed[3933],seed[470],seed[1148],seed[511],seed[586],seed[46],seed[1001],seed[631],seed[3162],seed[669],seed[1003],seed[2442],seed[2190],seed[3023],seed[3231],seed[261],seed[2083],seed[17],seed[3048],seed[812],seed[136],seed[3708],seed[1406],seed[390],seed[3877],seed[3823],seed[2653],seed[270],seed[958],seed[936],seed[1116],seed[2789],seed[2754],seed[1372],seed[164],seed[1264],seed[2385],seed[3952],seed[1731],seed[1978],seed[636],seed[397],seed[3640],seed[2944],seed[3199],seed[956],seed[1545],seed[1815],seed[1601],seed[3221],seed[2456],seed[1172],seed[1958],seed[3317],seed[2045],seed[1891],seed[2750],seed[3235],seed[3956],seed[39],seed[765],seed[2662],seed[2123],seed[1334],seed[45],seed[3695],seed[2271],seed[889],seed[3242],seed[2194],seed[3167],seed[1531],seed[2046],seed[1536],seed[3698],seed[2302],seed[3466],seed[3550],seed[2362],seed[2220],seed[1783],seed[249],seed[1962],seed[278],seed[930],seed[1035],seed[791],seed[929],seed[1796],seed[3248],seed[2966],seed[2634],seed[2455],seed[795],seed[2785],seed[3934],seed[1290],seed[1011],seed[1491],seed[3598],seed[2411],seed[425],seed[1275],seed[1008],seed[1801],seed[228],seed[284],seed[1774],seed[1251],seed[1305],seed[655],seed[1956],seed[2098],seed[1856],seed[2360],seed[4092],seed[3424],seed[2805],seed[1914],seed[3326],seed[2659],seed[4062],seed[1689],seed[1434],seed[412],seed[2576],seed[2586],seed[1664],seed[1030],seed[1982],seed[3145],seed[3100],seed[935],seed[622],seed[2751],seed[3440],seed[2877],seed[517],seed[419],seed[1896],seed[2610],seed[1379],seed[1260],seed[3484],seed[3007],seed[3959],seed[333],seed[2975],seed[3258],seed[1992],seed[1651],seed[1505],seed[497],seed[2612],seed[3862],seed[430],seed[2347],seed[1204],seed[3291],seed[3816],seed[1493],seed[141],seed[3212],seed[2429],seed[1947],seed[2682],seed[3376],seed[3509],seed[2386],seed[989],seed[321],seed[3965],seed[2809],seed[1794],seed[1199],seed[2737],seed[2939],seed[3335],seed[858],seed[1683],seed[778],seed[3252],seed[429],seed[1775],seed[768],seed[499],seed[3850],seed[3469],seed[2368],seed[632],seed[2249],seed[3652],seed[3519],seed[2334],seed[3285],seed[3473],seed[1534],seed[3375],seed[727],seed[1422],seed[111],seed[1843],seed[1122],seed[1424],seed[3264],seed[1750],seed[1441],seed[3441],seed[211],seed[2708],seed[3432],seed[2493],seed[3163],seed[1431],seed[1304],seed[1599],seed[759],seed[1705],seed[3430],seed[2930],seed[2649],seed[336],seed[2253],seed[590],seed[1739],seed[1259],seed[2824],seed[2047],seed[2650],seed[3800],seed[1282],seed[595],seed[2229],seed[810],seed[2890],seed[2434],seed[216],seed[1547],seed[2241],seed[475],seed[2257],seed[3233],seed[856],seed[2765],seed[494],seed[1912],seed[217],seed[1082],seed[2707],seed[1885],seed[1592],seed[2490],seed[1412],seed[2139],seed[965],seed[630],seed[3358],seed[1054],seed[245],seed[955],seed[451],seed[2954],seed[933],seed[4004],seed[2075],seed[4045],seed[149],seed[2683],seed[4053],seed[138],seed[2732],seed[2753],seed[1019],seed[4066],seed[644],seed[2248],seed[3052],seed[3896],seed[3147],seed[1697],seed[850],seed[297],seed[505],seed[60],seed[1127],seed[3569],seed[2672],seed[123],seed[1873],seed[2563],seed[2846],seed[4019],seed[839],seed[2461],seed[1691],seed[2444],seed[1711],seed[364],seed[373],seed[2950],seed[805],seed[3522],seed[2566],seed[1073],seed[1463],seed[1229],seed[1297],seed[2161],seed[1798],seed[4029],seed[3885],seed[1516],seed[1548],seed[3263],seed[606],seed[716],seed[3323],seed[3597],seed[3304],seed[251],seed[1614],seed[510],seed[2396],seed[3784],seed[1045],seed[1744],seed[3578],seed[1700],seed[2018],seed[3513],seed[4085],seed[90],seed[215],seed[365],seed[1039],seed[2121],seed[3299],seed[694],seed[2814],seed[2922],seed[1569],seed[1157],seed[1375],seed[773],seed[302],seed[2076],seed[1416],seed[2306],seed[3720],seed[1453],seed[2756],seed[1284],seed[1101],seed[3015],seed[140],seed[1849],seed[1460],seed[2114],seed[354],seed[1804],seed[377],seed[1155],seed[1507],seed[2230],seed[2397],seed[744],seed[3972],seed[2545],seed[1017],seed[1322],seed[3916],seed[659],seed[351],seed[104],seed[923],seed[3296],seed[4061],seed[2548],seed[2449],seed[137],seed[79],seed[1477],seed[798],seed[1524],seed[2092],seed[1608],seed[1378],seed[1443],seed[1826],seed[806],seed[1474],seed[2840],seed[3872],seed[452],seed[3731],seed[1254],seed[3680],seed[1778],seed[2422],seed[178],seed[641],seed[3058],seed[1440],seed[2870],seed[2131],seed[3420],seed[2579],seed[1139],seed[160],seed[1235],seed[3863],seed[2987],seed[712],seed[1883],seed[1456],seed[3261],seed[1971],seed[503],seed[4018],seed[3924],seed[3283],seed[561],seed[700],seed[3528],seed[2061],seed[1438],seed[2501],seed[241],seed[163],seed[1021],seed[3042],seed[1957],seed[2011],seed[3889],seed[2802],seed[1129],seed[2865],seed[2005],seed[1432],seed[3173],seed[2584],seed[3448],seed[2400],seed[789],seed[2670],seed[1317],seed[2568],seed[1162],seed[2286],seed[1294],seed[3943],seed[2729],seed[1863],seed[318],seed[2777],seed[1995],seed[2140],seed[1000],seed[2099],seed[1494],seed[2117],seed[2656],seed[786],seed[3101],seed[58],seed[2643],seed[2304],seed[3451],seed[36],seed[573],seed[3853],seed[1186],seed[3848],seed[3808],seed[1698],seed[3319],seed[2702],seed[3414],seed[3595],seed[1760],seed[2908],seed[4038],seed[3150],seed[2101],seed[2976],seed[3902],seed[2620],seed[3839],seed[1526],seed[2874],seed[2565],seed[3091],seed[482],seed[1185],seed[1837],seed[758],seed[2210],seed[1009],seed[1256],seed[781],seed[1280],seed[3325],seed[483],seed[1306],seed[4063],seed[3193],seed[1728],seed[3210],seed[571],seed[2658],seed[108],seed[2023],seed[3175],seed[645],seed[2948],seed[1184],seed[2974],seed[1944],seed[1435],seed[1931],seed[3401],seed[3754],seed[3805],seed[3761],seed[1541],seed[500],seed[1542],seed[2989],seed[591],seed[717],seed[2425],seed[4088],seed[3211],seed[1024],seed[421],seed[1661],seed[2710],seed[348],seed[3392],seed[612],seed[1951],seed[2627],seed[15],seed[1701],seed[3904],seed[2760],seed[2863],seed[1403],seed[1954],seed[704],seed[3579],seed[2291],seed[3673],seed[2015],seed[3886],seed[1156],seed[3382],seed[2641],seed[2764],seed[803],seed[3017],seed[1038],seed[3922],seed[3810],seed[461],seed[3179],seed[629],seed[589],seed[1223],seed[2149],seed[2781],seed[2152],seed[3832],seed[2082],seed[1452],seed[2907],seed[1656],seed[943],seed[3964],seed[1650],seed[446],seed[1824],seed[1588],seed[197],seed[1158],seed[3549],seed[2958],seed[512],seed[3228],seed[3236],seed[1960],seed[4020],seed[350],seed[2084],seed[1094],seed[1842],seed[829],seed[1964],seed[189],seed[3316],seed[1049],seed[3348],seed[1573],seed[619],seed[3606],seed[2293],seed[188],seed[1718],seed[2704],seed[3246],seed[3767],seed[3185],seed[382],seed[1765],seed[1271],seed[3201],seed[1108],seed[3064],seed[2193],seed[2798],seed[346],seed[1149],seed[973],seed[3676],seed[2314],seed[2470],seed[1272],seed[2716],seed[2847],seed[2577],seed[122],seed[33],seed[992],seed[3925],seed[1263],seed[1764],seed[525],seed[2744],seed[3388],seed[3374],seed[2219],seed[2124],seed[807],seed[247],seed[1763],seed[1091],seed[1519],seed[471],seed[702],seed[3892],seed[3947],seed[4046],seed[3537],seed[2538],seed[2766],seed[116],seed[1490],seed[3693],seed[1346],seed[78],seed[2995],seed[3530],seed[2031],seed[2736],seed[2127],seed[2315],seed[239],seed[3284],seed[502],seed[82],seed[3529],seed[176],seed[3748],seed[1083],seed[1439],seed[2182],seed[677],seed[838],seed[2159],seed[320],seed[3732],seed[1979],seed[1351],seed[3391],seed[3226],seed[551],seed[1340],seed[1632],seed[2361],seed[4044],seed[3313],seed[2421],seed[2504],seed[2327],seed[4079],seed[2441],seed[667],seed[3407],seed[3223],seed[2469],seed[363],seed[225],seed[3144],seed[835],seed[1090],seed[3700],seed[897],seed[3485],seed[1732],seed[2478],seed[3931],seed[1338],seed[2875],seed[3681],seed[1754],seed[2558],seed[1867],seed[1868],seed[3217],seed[3527],seed[2192],seed[324],seed[1727],seed[2723],seed[2832],seed[1196],seed[2990],seed[14],seed[1471],seed[2363],seed[3604],seed[2943],seed[2884],seed[3218],seed[860],seed[1060],seed[890],seed[2198],seed[26],seed[3600],seed[1010],seed[642],seed[1245],seed[1512],seed[2748],seed[4041],seed[4000],seed[1448],seed[1864],seed[3704],seed[6],seed[736],seed[3768],seed[711],seed[2108],seed[3396],seed[2921],seed[2506],seed[3403],seed[2086],seed[2336],seed[1190],seed[1981],seed[2435],seed[3125],seed[1119],seed[2703],seed[1472],seed[3814],seed[2163],seed[1459],seed[3987],seed[3524],seed[1429],seed[513],seed[2984],seed[1915],seed[47],seed[1603],seed[1594],seed[1145],seed[3498],seed[1087],seed[238],seed[3307],seed[424],seed[1670],seed[3894],seed[3416],seed[3584],seed[2164],seed[2836],seed[1695],seed[687],seed[3697],seed[2231],seed[2319],seed[2735],seed[3562],seed[465],seed[721],seed[69],seed[4072],seed[1323],seed[1630],seed[3900],seed[349],seed[3080],seed[2848],seed[847],seed[2172],seed[3131],seed[76],seed[3274],seed[3914],seed[98],seed[1257],seed[1426],seed[3817],seed[307],seed[766],seed[2618],seed[556],seed[3298],seed[1068],seed[19],seed[699],seed[2473],seed[2691],seed[2539],seed[1974],seed[148],seed[2016],seed[2338],seed[481],seed[3337],seed[1164],seed[1207],seed[3450],seed[303],seed[2556],seed[2537],seed[3072],seed[132],seed[865],seed[366],seed[902],seed[1369],seed[3594],seed[726],seed[3646],seed[2268],seed[1262],seed[2285],seed[269],seed[1851],seed[1138],seed[1401],seed[2142],seed[396],seed[1741],seed[3560],seed[1539],seed[367],seed[1299],seed[308],seed[817],seed[594],seed[1919],seed[1803],seed[3096],seed[1075],seed[2070],seed[3857],seed[2685],seed[3279],seed[2356],seed[3670],seed[2999],seed[1012],seed[2878],seed[3561],seed[975],seed[605],seed[1602],seed[3419],seed[3196],seed[89],seed[3899],seed[300],seed[3437],seed[1517],seed[3390],seed[1621],seed[355],seed[3706],seed[637],seed[1570],seed[2792],seed[3355],seed[2779],seed[370],seed[454],seed[53],seed[3363],seed[3204],seed[3427],seed[725],seed[3483],seed[1777],seed[2550],seed[2714],seed[2902],seed[2889],seed[1048],seed[2322],seed[1871],seed[1955],seed[2869],seed[2853],seed[2740],seed[3362],seed[3514],seed[2800],seed[1953],seed[1950],seed[1215],seed[906],seed[609],seed[3559],seed[456],seed[3614],seed[3068],seed[2898],seed[649],seed[3132],seed[964],seed[3053],seed[1899],seed[220],seed[2582],seed[508],seed[1309],seed[2838],seed[535],seed[2615],seed[329],seed[177],seed[1395],seed[2739],seed[3057],seed[119],seed[1007],seed[522],seed[3912],seed[2038],seed[1716],seed[3735],seed[3310],seed[2823],seed[756],seed[4027],seed[2367],seed[4084],seed[1026],seed[473],seed[809],seed[3000],seed[2333],seed[1462],seed[1399],seed[1480],seed[1903],seed[1407],seed[993],seed[337],seed[962],seed[2081],seed[3148],seed[1069],seed[802],seed[2619],seed[2589],seed[2856],seed[2433],seed[2928],seed[2813],seed[2175],seed[1706],seed[1391],seed[743],seed[327],seed[1345],seed[1677],seed[2032],seed[394],seed[3994],seed[3861],seed[4014],seed[1197],seed[899],seed[3453],seed[1332],seed[1787],seed[2758],seed[3275],seed[3723],seed[3143],seed[1250],seed[194],seed[4058],seed[3884],seed[28],seed[1527],seed[1253],seed[3339],seed[904],seed[2978],seed[3288],seed[1707],seed[2852],seed[1736],seed[2317],seed[3151],seed[3874],seed[514],seed[3954],seed[1726],seed[1942],seed[3826],seed[361],seed[2165],seed[1377],seed[345],seed[2894],seed[1454],seed[3181],seed[1002],seed[831],seed[3710],seed[1444],seed[1788],seed[3454],seed[2244],seed[826],seed[3517],seed[1201],seed[757],seed[3938],seed[1059],seed[3962],seed[2111],seed[50],seed[1086],seed[3669],seed[2912],seed[3541],seed[2859],seed[568],seed[2450],seed[2453],seed[915],seed[731],seed[1140],seed[2951],seed[444],seed[921],seed[945],seed[1469],seed[2913],seed[10],seed[2122],seed[2699],seed[1789],seed[3953],seed[578],seed[1041],seed[356],seed[967],seed[3993],seed[2614],seed[2666],seed[800],seed[2072],seed[2062],seed[1504],seed[1034],seed[2344],seed[2742],seed[165],seed[2745],seed[3539],seed[1595],seed[3613],seed[608],seed[1133],seed[1638],seed[1072],seed[2498],seed[32],seed[1666],seed[521],seed[1478],seed[1110],seed[2988],seed[3782],seed[3687],seed[2412],seed[604],seed[1052],seed[1756],seed[3146],seed[314],seed[3063],seed[2048],seed[3043],seed[3821],seed[2596],seed[4073],seed[912],seed[443],seed[536],seed[3905],seed[3215],seed[191],seed[2561],seed[2189],seed[190],seed[3656],seed[2406],seed[2346],seed[3563],seed[3834],seed[3230],seed[2717],seed[2973],seed[4013],seed[2339],seed[1370],seed[3958],seed[2144],seed[868],seed[1291],seed[3489],seed[74],seed[1772],seed[2279],seed[5],seed[4076],seed[584],seed[2552],seed[3664],seed[2395],seed[2505],seed[1563],seed[31],seed[3379],seed[3036],seed[2960],seed[914],seed[1099],seed[3014],seed[1965],seed[3713],seed[729],seed[3622],seed[3314],seed[748],seed[1449],seed[3384],seed[2151],seed[3495],seed[2486],seed[2830],seed[1721],seed[3996],seed[3675],seed[3696],seed[3031],seed[1043],seed[3567],seed[3980],seed[1225],seed[1712],seed[4003],seed[1255],seed[3984],seed[3608],seed[1065],seed[724],seed[1799],seed[1874],seed[3084],seed[1847],seed[2786],seed[2844],seed[683],seed[3534],seed[949],seed[3688],seed[698],seed[2495],seed[3525],seed[3571],seed[3281],seed[476],seed[3715],seed[601],seed[919],seed[387],seed[2808],seed[2711],seed[323],seed[48],seed[549],seed[1163],seed[544],seed[3460],seed[1671],seed[3751],seed[273],seed[3174],seed[401],seed[3662],seed[408],seed[3679],seed[2799],seed[3729],seed[652]};
//        seed2 <= {seed[3755],seed[988],seed[3960],seed[2859],seed[2044],seed[1829],seed[2116],seed[1015],seed[1573],seed[1704],seed[2775],seed[3485],seed[652],seed[3089],seed[3870],seed[2905],seed[697],seed[1077],seed[1635],seed[2457],seed[1786],seed[337],seed[2174],seed[101],seed[2450],seed[3605],seed[2850],seed[2035],seed[2159],seed[3982],seed[1114],seed[3291],seed[3289],seed[3535],seed[1626],seed[1554],seed[853],seed[748],seed[1319],seed[1394],seed[3878],seed[2749],seed[689],seed[129],seed[1527],seed[3544],seed[590],seed[1489],seed[3025],seed[3055],seed[187],seed[3351],seed[744],seed[814],seed[507],seed[1270],seed[2474],seed[2639],seed[2600],seed[1353],seed[2841],seed[598],seed[3751],seed[1558],seed[3747],seed[1323],seed[746],seed[1875],seed[2814],seed[800],seed[4054],seed[1390],seed[180],seed[3702],seed[1134],seed[1138],seed[761],seed[874],seed[3410],seed[3995],seed[3958],seed[416],seed[4061],seed[3700],seed[585],seed[1706],seed[2538],seed[733],seed[2874],seed[1736],seed[449],seed[985],seed[2307],seed[54],seed[1898],seed[712],seed[3431],seed[856],seed[150],seed[727],seed[1537],seed[774],seed[1305],seed[2867],seed[2722],seed[721],seed[2616],seed[1284],seed[2017],seed[1456],seed[68],seed[2106],seed[4089],seed[3593],seed[1686],seed[364],seed[208],seed[2570],seed[919],seed[1940],seed[3326],seed[1079],seed[880],seed[3484],seed[961],seed[3411],seed[2279],seed[495],seed[888],seed[1807],seed[3013],seed[2382],seed[1619],seed[2120],seed[1004],seed[1980],seed[2950],seed[1605],seed[297],seed[2322],seed[3518],seed[1989],seed[1910],seed[1580],seed[2014],seed[1225],seed[1974],seed[506],seed[1876],seed[3557],seed[3369],seed[3546],seed[1363],seed[3770],seed[4035],seed[2624],seed[2271],seed[3576],seed[3930],seed[665],seed[1239],seed[3395],seed[3111],seed[3365],seed[3635],seed[2986],seed[3421],seed[3831],seed[2376],seed[312],seed[1998],seed[1287],seed[3683],seed[1852],seed[1480],seed[661],seed[1691],seed[3618],seed[1006],seed[3667],seed[2261],seed[4030],seed[1497],seed[244],seed[340],seed[3904],seed[3820],seed[2419],seed[1911],seed[1777],seed[3743],seed[1314],seed[3956],seed[3312],seed[1016],seed[350],seed[1375],seed[1117],seed[3246],seed[3631],seed[2893],seed[1423],seed[3415],seed[2422],seed[39],seed[3465],seed[3414],seed[1279],seed[2223],seed[2292],seed[2621],seed[3451],seed[3556],seed[3693],seed[1013],seed[1962],seed[3745],seed[715],seed[618],seed[3496],seed[3974],seed[2987],seed[3838],seed[2999],seed[3200],seed[3052],seed[140],seed[1514],seed[1630],seed[2104],seed[351],seed[4057],seed[4060],seed[2585],seed[1106],seed[3458],seed[1121],seed[957],seed[3595],seed[3638],seed[2448],seed[964],seed[656],seed[1377],seed[1078],seed[863],seed[1740],seed[2804],seed[1281],seed[2820],seed[2612],seed[807],seed[1617],seed[3011],seed[1871],seed[1930],seed[1470],seed[2752],seed[3066],seed[3021],seed[1963],seed[3905],seed[3777],seed[2015],seed[605],seed[1830],seed[2598],seed[2653],seed[1792],seed[135],seed[2484],seed[829],seed[2695],seed[1419],seed[2383],seed[2206],seed[3876],seed[430],seed[182],seed[3252],seed[1739],seed[3007],seed[1929],seed[250],seed[1559],seed[1782],seed[367],seed[594],seed[2565],seed[1757],seed[629],seed[1781],seed[824],seed[3785],seed[3815],seed[3215],seed[846],seed[3714],seed[927],seed[305],seed[3146],seed[2561],seed[3071],seed[3599],seed[4049],seed[3880],seed[3294],seed[3726],seed[1943],seed[3076],seed[553],seed[3059],seed[1009],seed[2700],seed[510],seed[2034],seed[2471],seed[59],seed[3773],seed[2916],seed[959],seed[2493],seed[749],seed[3727],seed[418],seed[282],seed[546],seed[262],seed[3340],seed[96],seed[3711],seed[338],seed[2674],seed[2951],seed[539],seed[3148],seed[3017],seed[693],seed[3607],seed[429],seed[2808],seed[2053],seed[840],seed[3302],seed[1436],seed[1841],seed[1324],seed[986],seed[1112],seed[319],seed[138],seed[3429],seed[3695],seed[516],seed[3149],seed[3166],seed[2851],seed[706],seed[1195],seed[2529],seed[4083],seed[2932],seed[1049],seed[222],seed[384],seed[163],seed[2890],seed[2815],seed[969],seed[1799],seed[291],seed[3975],seed[2954],seed[1442],seed[2944],seed[34],seed[467],seed[3152],seed[3416],seed[3924],seed[531],seed[3268],seed[2679],seed[4062],seed[1250],seed[595],seed[675],seed[153],seed[1310],seed[2738],seed[3664],seed[2568],seed[315],seed[2154],seed[2233],seed[2756],seed[3676],seed[1627],seed[3879],seed[520],seed[3996],seed[3644],seed[236],seed[2992],seed[1027],seed[2998],seed[1298],seed[2548],seed[827],seed[1268],seed[1304],seed[1983],seed[869],seed[3571],seed[2761],seed[809],seed[2193],seed[69],seed[3792],seed[3186],seed[698],seed[3629],seed[2681],seed[162],seed[3944],seed[1482],seed[3718],seed[2983],seed[2685],seed[1730],seed[3028],seed[3784],seed[1376],seed[1414],seed[1770],seed[2648],seed[1572],seed[597],seed[3740],seed[2298],seed[3673],seed[3603],seed[2521],seed[3843],seed[3407],seed[1759],seed[46],seed[2751],seed[2147],seed[1897],seed[2978],seed[3437],seed[448],seed[2153],seed[2100],seed[1160],seed[1382],seed[2614],seed[3251],seed[3277],seed[3990],seed[3135],seed[601],seed[1251],seed[617],seed[789],seed[1211],seed[4050],seed[716],seed[2296],seed[2184],seed[3347],seed[2288],seed[3889],seed[4064],seed[730],seed[207],seed[486],seed[1564],seed[555],seed[1407],seed[155],seed[1976],seed[682],seed[2675],seed[1655],seed[3621],seed[1206],seed[491],seed[3453],seed[3789],seed[1005],seed[3528],seed[2750],seed[261],seed[1043],seed[3232],seed[1970],seed[3947],seed[2370],seed[2941],seed[333],seed[1519],seed[1510],seed[3156],seed[2563],seed[1848],seed[1269],seed[947],seed[3907],seed[902],seed[3931],seed[509],seed[2929],seed[778],seed[1296],seed[1701],seed[2901],seed[982],seed[3202],seed[2152],seed[1902],seed[198],seed[2062],seed[2844],seed[2140],seed[3520],seed[3688],seed[784],seed[2308],seed[3053],seed[382],seed[1431],seed[2723],seed[1529],seed[1997],seed[3479],seed[183],seed[2619],seed[3509],seed[723],seed[1645],seed[1007],seed[1194],seed[1168],seed[2086],seed[308],seed[1889],seed[341],seed[2222],seed[2213],seed[1430],seed[780],seed[1666],seed[3412],seed[3067],seed[1209],seed[3766],seed[662],seed[3385],seed[1958],seed[492],seed[695],seed[1561],seed[1397],seed[1371],seed[1754],seed[108],seed[424],seed[604],seed[2762],seed[2402],seed[3712],seed[3138],seed[1637],seed[175],seed[900],seed[4004],seed[2584],seed[2314],seed[1062],seed[1399],seed[293],seed[2914],seed[2161],seed[3886],seed[980],seed[3370],seed[4065],seed[1245],seed[158],seed[521],seed[130],seed[2212],seed[1110],seed[3307],seed[3682],seed[3660],seed[2855],seed[254],seed[2609],seed[9],seed[2937],seed[3454],seed[2861],seed[3636],seed[758],seed[511],seed[3519],seed[527],seed[422],seed[1339],seed[573],seed[2395],seed[299],seed[2165],seed[3853],seed[3567],seed[3937],seed[1347],seed[3661],seed[389],seed[3267],seed[2096],seed[1815],seed[1498],seed[2650],seed[794],seed[3387],seed[3271],seed[3882],seed[1813],seed[2627],seed[2657],seed[3086],seed[2838],seed[2730],seed[2210],seed[3494],seed[1299],seed[1357],seed[202],seed[322],seed[420],seed[2134],seed[2012],seed[3273],seed[1349],seed[2965],seed[51],seed[2935],seed[74],seed[967],seed[1212],seed[3457],seed[2172],seed[1023],seed[1745],seed[2342],seed[1996],seed[2879],seed[3901],seed[2185],seed[154],seed[85],seed[3078],seed[2214],seed[215],seed[3570],seed[2728],seed[1530],seed[2175],seed[1122],seed[3809],seed[1396],seed[3476],seed[2257],seed[3652],seed[1622],seed[848],seed[1180],seed[3339],seed[1022],seed[2275],seed[3912],seed[1141],seed[2158],seed[2238],seed[289],seed[2355],seed[569],seed[3217],seed[3506],seed[1649],seed[565],seed[2871],seed[1142],seed[1845],seed[2490],seed[2235],seed[1364],seed[1668],seed[2125],seed[2323],seed[3213],seed[1085],seed[3617],seed[318],seed[994],seed[230],seed[3909],seed[2516],seed[2114],seed[415],seed[632],seed[909],seed[951],seed[1317],seed[1964],seed[2203],seed[649],seed[645],seed[1948],seed[1176],seed[3706],seed[1583],seed[1352],seed[3609],seed[1960],seed[3753],seed[1609],seed[2806],seed[3128],seed[460],seed[4042],seed[3736],seed[953],seed[2899],seed[3869],seed[2121],seed[219],seed[1385],seed[3994],seed[103],seed[1837],seed[88],seed[885],seed[3503],seed[2766],seed[3633],seed[4071],seed[410],seed[2888],seed[2961],seed[157],seed[567],seed[2290],seed[523],seed[3285],seed[641],seed[457],seed[160],seed[400],seed[223],seed[2434],seed[1586],seed[3689],seed[1779],seed[3101],seed[4017],seed[3493],seed[1593],seed[3950],seed[2705],seed[136],seed[2108],seed[2351],seed[786],seed[2072],seed[2956],seed[924],seed[3906],seed[2958],seed[1823],seed[2880],seed[2683],seed[1767],seed[2854],seed[3112],seed[2039],seed[1500],seed[2835],seed[271],seed[2091],seed[1766],seed[2664],seed[561],seed[2805],seed[3207],seed[530],seed[3619],seed[1624],seed[2302],seed[1097],seed[1629],seed[248],seed[19],seed[2892],seed[2803],seed[2549],seed[2135],seed[1053],seed[1320],seed[3548],seed[1291],seed[628],seed[1157],seed[3697],seed[2483],seed[1466],seed[2939],seed[3296],seed[1208],seed[816],seed[547],seed[1654],seed[177],seed[918],seed[2923],seed[2389],seed[996],seed[485],seed[732],seed[2727],seed[1746],seed[4095],seed[3471],seed[3835],seed[972],seed[3829],seed[1824],seed[529],seed[2863],seed[2515],seed[1453],seed[73],seed[394],seed[4053],seed[1771],seed[3513],seed[4015],seed[3206],seed[390],seed[1205],seed[3191],seed[3516],seed[253],seed[737],seed[3921],seed[2885],seed[1204],seed[2128],seed[2057],seed[2647],seed[2503],seed[3171],seed[3709],seed[2967],seed[2597],seed[3733],seed[1031],seed[680],seed[1484],seed[164],seed[2010],seed[3504],seed[3033],seed[2702],seed[3464],seed[440],seed[206],seed[971],seed[830],seed[575],seed[292],seed[2847],seed[1018],seed[993],seed[912],seed[592],seed[3338],seed[1661],seed[4067],seed[3978],seed[1667],seed[2966],seed[316],seed[3137],seed[3648],seed[4036],seed[89],seed[3314],seed[2478],seed[3642],seed[3678],seed[1086],seed[2712],seed[2295],seed[3438],seed[2862],seed[3954],seed[1330],seed[3258],seed[2240],seed[2348],seed[872],seed[1715],seed[1246],seed[2102],seed[1546],seed[3113],seed[1720],seed[52],seed[1452],seed[4052],seed[775],seed[2662],seed[3898],seed[1064],seed[210],seed[489],seed[1136],seed[2560],seed[3325],seed[1116],seed[311],seed[3490],seed[2004],seed[2332],seed[965],seed[2263],seed[3189],seed[2535],seed[1181],seed[2189],seed[1354],seed[3379],seed[2453],seed[3220],seed[2799],seed[2786],seed[1615],seed[2668],seed[2477],seed[1446],seed[487],seed[2949],seed[1955],seed[1461],seed[3797],seed[233],seed[2069],seed[2920],seed[2306],seed[1680],seed[2607],seed[3293],seed[2473],seed[2637],seed[2573],seed[3359],seed[3115],seed[3641],seed[570],seed[3272],seed[456],seed[2347],seed[709],seed[1153],seed[2593],seed[1838],seed[399],seed[3276],seed[2699],seed[1036],seed[3803],seed[2928],seed[8],seed[1381],seed[1095],seed[3545],seed[3175],seed[1513],seed[442],seed[3943],seed[2718],seed[3139],seed[2532],seed[3160],seed[781],seed[1081],seed[823],seed[2669],seed[958],seed[3009],seed[788],seed[3948],seed[1696],seed[2460],seed[1221],seed[1263],seed[704],seed[3914],seed[1731],seed[117],seed[3341],seed[1282],seed[3110],seed[1140],seed[3505],seed[228],seed[4058],seed[1589],seed[679],seed[1869],seed[1576],seed[2737],seed[2865],seed[2527],seed[3436],seed[423],seed[2789],seed[3245],seed[538],seed[3125],seed[3243],seed[1236],seed[519],seed[3036],seed[2747],seed[3897],seed[1984],seed[710],seed[1285],seed[3211],seed[2782],seed[2426],seed[2580],seed[1014],seed[4045],seed[1459],seed[837],seed[124],seed[1679],seed[331],seed[3116],seed[1550],seed[822],seed[1538],seed[2623],seed[2058],seed[3507],seed[344],seed[3363],seed[1855],seed[25],seed[3888],seed[3153],seed[3380],seed[3925],seed[4007],seed[1517],seed[3345],seed[1785],seed[542],seed[417],seed[3604],seed[3157],seed[76],seed[3499],seed[1863],seed[13],seed[633],seed[1473],seed[2542],seed[67],seed[1728],seed[1856],seed[2216],seed[3404],seed[329],seed[1947],seed[2595],seed[335],seed[1794],seed[2231],seed[1692],seed[1093],seed[2280],seed[1108],seed[1173],seed[1651],seed[1326],seed[1297],seed[771],seed[3971],seed[143],seed[883],seed[3854],seed[2823],seed[1698],seed[1019],seed[2821],seed[502],seed[3615],seed[2377],seed[2282],seed[4000],seed[3440],seed[476],seed[2368],seed[3095],seed[2007],seed[1543],seed[243],seed[3722],seed[2895],seed[403],seed[3281],seed[1893],seed[3366],seed[3981],seed[3832],seed[225],seed[4023],seed[3495],seed[2707],seed[847],seed[2617],seed[3234],seed[60],seed[2971],seed[990],seed[1230],seed[2437],seed[2363],seed[3039],seed[4076],seed[4019],seed[113],seed[747],seed[2759],seed[640],seed[1542],seed[3424],seed[1226],seed[941],seed[3614],seed[3685],seed[1750],seed[893],seed[3342],seed[1697],seed[2973],seed[2379],seed[2466],seed[4027],seed[2499],seed[239],seed[104],seed[2903],seed[234],seed[2482],seed[1045],seed[1791],seed[1432],seed[1709],seed[3561],seed[1532],seed[700],seed[2463],seed[2725],seed[4094],seed[365],seed[2136],seed[2447],seed[285],seed[2469],seed[669],seed[2876],seed[1826],seed[745],seed[3330],seed[862],seed[378],seed[1096],seed[1986],seed[1469],seed[1336],seed[3391],seed[678],seed[4006],seed[2180],seed[3131],seed[200],seed[2415],seed[1101],seed[452],seed[1126],seed[841],seed[2846],seed[1415],seed[696],seed[1207],seed[2760],seed[2160],seed[310],seed[4056],seed[1999],seed[798],seed[1858],seed[357],seed[3526],seed[1665],seed[1919],seed[634],seed[3515],seed[2663],seed[3237],seed[648],seed[2975],seed[1272],seed[3775],seed[224],seed[2250],seed[1507],seed[4003],seed[1425],seed[3899],seed[1951],seed[3840],seed[2051],seed[2101],seed[3389],seed[2801],seed[3275],seed[1935],seed[2429],seed[549],seed[2922],seed[1198],seed[2038],seed[2026],seed[1197],seed[4010],seed[82],seed[690],seed[77],seed[435],seed[2470],seed[3579],seed[1408],seed[2673],seed[3744],seed[1429],seed[2770],seed[3127],seed[2398],seed[677],seed[2646],seed[1151],seed[3824],seed[36],seed[4079],seed[1312],seed[2601],seed[2391],seed[624],seed[336],seed[2656],seed[3554],seed[1660],seed[2860],seed[106],seed[3560],seed[708],seed[2566],seed[2757],seed[3798],seed[120],seed[3238],seed[2365],seed[3502],seed[3032],seed[2050],seed[3332],seed[3195],seed[2107],seed[2392],seed[2090],seed[23],seed[184],seed[3406],seed[1894],seed[1805],seed[3932],seed[3764],seed[2710],seed[1836],seed[2232],seed[275],seed[3668],seed[2740],seed[1941],seed[3591],seed[861],seed[540],seed[231],seed[3517],seed[4082],seed[2186],seed[1975],seed[3483],seed[3107],seed[1934],seed[916],seed[1844],seed[201],seed[2319],seed[3382],seed[884],seed[3320],seed[3872],seed[105],seed[2817],seed[3836],seed[2583],seed[2412],seed[1772],seed[831],seed[141],seed[3821],seed[1670],seed[3018],seed[2143],seed[1891],seed[2028],seed[1069],seed[3123],seed[2955],seed[1909],seed[3247],seed[2701],seed[2046],seed[4016],seed[2825],seed[1169],seed[1188],seed[3655],seed[797],seed[2179],seed[2061],seed[2413],seed[3555],seed[3208],seed[220],seed[3696],seed[929],seed[4048],seed[688],seed[251],seed[2097],seed[4033],seed[1384],seed[1795],seed[2495],seed[1174],seed[3260],seed[1928],seed[3420],seed[1783],seed[65],seed[2795],seed[2665],seed[3224],seed[2094],seed[1088],seed[528],seed[1398],seed[3169],seed[2582],seed[1601],seed[3558],seed[3178],seed[1927],seed[1711],seed[1274],seed[843],seed[3346],seed[1041],seed[579],seed[804],seed[2635],seed[1907],seed[2845],seed[653],seed[3527],seed[2224],seed[3003],seed[599],seed[466],seed[937],seed[3769],seed[1026],seed[2278],seed[1872],seed[2947],seed[3394],seed[1133],seed[2171],seed[431],seed[2170],seed[3933],seed[3060],seed[1575],seed[583],seed[375],seed[404],seed[3691],seed[956],seed[2887],seed[2373],seed[407],seed[3073],seed[2514],seed[332],seed[3934],seed[49],seed[266],seed[2011],seed[3825],seed[821],seed[1784],seed[3540],seed[718],seed[2401],seed[2792],seed[342],seed[1659],seed[1039],seed[1954],seed[369],seed[3396],seed[3158],seed[3108],seed[1977],seed[12],seed[3757],seed[891],seed[3235],seed[805],seed[2918],seed[1061],seed[2643],seed[672],seed[811],seed[3362],seed[1420],seed[286],seed[212],seed[2993],seed[1258],seed[955],seed[465],seed[3525],seed[2713],seed[844],seed[3857],seed[1071],seed[1146],seed[1387],seed[2076],seed[2872],seed[808],seed[1877],seed[3827],seed[2571],seed[3063],seed[392],seed[2547],seed[4088],seed[2997],seed[2802],seed[196],seed[1663],seed[3057],seed[3430],seed[3720],seed[40],seed[3632],seed[3628],seed[1228],seed[2852],seed[3000],seed[666],seed[1224],seed[1641],seed[2704],seed[3596],seed[515],seed[3304],seed[2192],seed[2071],seed[2324],seed[2018],seed[3481],seed[3855],seed[413],seed[2940],seed[2843],seed[4032],seed[1604],seed[2790],seed[55],seed[1918],seed[1454],seed[2708],seed[3222],seed[3278],seed[548],seed[1683],seed[371],seed[4063],seed[1],seed[1677],seed[1717],seed[2080],seed[3608],seed[2896],seed[2145],seed[2444],seed[3368],seed[2118],seed[623],seed[3957],seed[1778],seed[1074],seed[3223],seed[3069],seed[3936],seed[921],seed[21],seed[1293],seed[2113],seed[3928],seed[2518],seed[2869],seed[3643],seed[1082],seed[2042],seed[881],seed[2558],seed[482],seed[2574],seed[1578],seed[2645],seed[1551],seed[1648],seed[724],seed[139],seed[3480],seed[2191],seed[3445],seed[533],seed[2731],seed[3257],seed[612],seed[1994],seed[2139],seed[731],seed[3002],seed[2253],seed[2181],seed[2743],seed[796],seed[550],seed[3197],seed[740],seed[1913],seed[2546],seed[1276],seed[2837],seed[987],seed[536],seed[759],seed[1424],seed[144],seed[770],seed[169],seed[2268],seed[453],seed[2411],seed[2251],seed[3622],seed[43],seed[2606],seed[932],seed[2047],seed[3261],seed[1761],seed[588],seed[1985],seed[580],seed[2906],seed[3219],seed[2227],seed[1887],seed[2052],seed[2716],seed[1137],seed[2099],seed[2427],seed[3626],seed[4008],seed[1528],seed[2040],seed[3795],seed[908],seed[1524],seed[1266],seed[2089],seed[3162],seed[2828],seed[806],seed[2449],seed[2926],seed[1652],seed[112],seed[2375],seed[1865],seed[3814],seed[2894],seed[674],seed[2310],seed[1159],seed[2327],seed[2996],seed[3765],seed[735],seed[3724],seed[1467],seed[1416],seed[2953],seed[3731],seed[1154],seed[3637],seed[2221],seed[3917],seed[743],seed[2959],seed[2649],seed[1494],seed[3601],seed[3180],seed[2423],seed[2334],seed[767],seed[2618],seed[850],seed[1201],seed[1118],seed[3521],seed[1373],seed[2273],seed[3274],seed[1705],seed[1850],seed[564],seed[2689],seed[3910],seed[3828],seed[1802],seed[3951],seed[115],seed[147],seed[1769],seed[3375],seed[3598],seed[4005],seed[3692],seed[1688],seed[2019],seed[1816],seed[2318],seed[3093],seed[114],seed[1318],seed[3704],seed[2505],seed[3042],seed[3799],seed[1890],seed[3998],seed[1541],seed[3987],seed[2900],seed[2380],seed[2672],seed[2151],seed[2839],seed[3826],seed[1922],seed[3877],seed[127],seed[1789],seed[1614],seed[3164],seed[2556],seed[2927],seed[657],seed[2367],seed[81],seed[3543],seed[3941],seed[3145],seed[324],seed[4068],seed[1669],seed[3589],seed[501],seed[2305],seed[1215],seed[2182],seed[2098],seed[178],seed[2496],seed[2487],seed[4092],seed[2024],seed[2698],seed[1516],seed[2283],seed[2265],seed[2753],seed[2336],seed[1574],seed[2311],seed[545],seed[4046],seed[1451],seed[2462],seed[1884],seed[2857],seed[3707],seed[1846],seed[3865],seed[3462],seed[170],seed[1747],seed[3126],seed[1582],seed[1762],seed[673],seed[952],seed[1441],seed[111],seed[3737],seed[80],seed[2919],seed[2127],seed[2576],seed[6],seed[1072],seed[1010],seed[3913],seed[946],seed[2043],seed[2729],seed[277],seed[2122],seed[1867],seed[3742],seed[205],seed[84],seed[3225],seed[685],seed[1639],seed[3097],seed[2765],seed[1162],seed[216],seed[865],seed[358],seed[1623],seed[2141],seed[915],seed[2027],seed[877],seed[4039],seed[276],seed[2798],seed[1694],seed[295],seed[1506],seed[3204],seed[93],seed[2312],seed[2079],seed[2016],seed[2776],seed[398],seed[3360],seed[4072],seed[1793],seed[3241],seed[1636],seed[3012],seed[2432],seed[3734],seed[1981],seed[3647],seed[31],seed[1428],seed[832],seed[3199],seed[1926],seed[3443],seed[2316],seed[2533],seed[3315],seed[3151],seed[637],seed[3927],seed[734],seed[3068],seed[3659],seed[1040],seed[3967],seed[2344],seed[868],seed[1368],seed[3161],seed[1184],seed[896],seed[1650],seed[2651],seed[1565],seed[554],seed[833],seed[2162],seed[562],seed[572],seed[2048],seed[1768],seed[2671],seed[1389],seed[2946],seed[2281],seed[1075],seed[522],seed[1275],seed[3284],seed[1308],seed[1833],seed[1931],seed[1148],seed[2575],seed[3433],seed[3122],seed[907],seed[684],seed[541],seed[3300],seed[3035],seed[1254],seed[736],seed[2824],seed[1818],seed[2562],seed[374],seed[2301],seed[2372],seed[2758],seed[2544],seed[4020],seed[2362],seed[574],seed[3231],seed[2764],seed[3085],seed[1870],seed[875],seed[764],seed[1904],seed[1673],seed[566],seed[1400],seed[3719],seed[871],seed[2613],seed[1883],seed[1278],seed[193],seed[2693],seed[2243],seed[1952],seed[991],seed[2523],seed[4024],seed[2554],seed[2615],seed[1448],seed[2218],seed[934],seed[3045],seed[3102],seed[2706],seed[2060],seed[1812],seed[1046],seed[3552],seed[3333],seed[4025],seed[1147],seed[1625],seed[2994],seed[935],seed[2884],seed[1968],seed[2735],seed[857],seed[4040],seed[2970],seed[512],seed[3830],seed[1643],seed[2220],seed[211],seed[763],seed[3254],seed[2260],seed[2811],seed[2315],seed[3316],seed[984],seed[1238],seed[1163],seed[161],seed[2632],seed[2359],seed[1232],seed[1322],seed[107],seed[3027],seed[3542],seed[867],seed[499],seed[4051],seed[1503],seed[1288],seed[3962],seed[1050],seed[1035],seed[3323],seed[444],seed[1713],seed[2188],seed[3472],seed[2721],seed[1886],seed[1658],seed[3061],seed[1504],seed[596],seed[3079],seed[1840],seed[1161],seed[3313],seed[1068],seed[1348],seed[3966],seed[819],seed[1949],seed[4014],seed[1488],seed[1882],seed[1143],seed[3915],seed[2123],seed[1367],seed[2781],seed[370],seed[1776],seed[1827],seed[1773],seed[3781],seed[2769],seed[2777],seed[98],seed[2506],seed[2406],seed[2744],seed[1920],seed[1515],seed[438],seed[1612],seed[3823],seed[1721],seed[1025],seed[2196],seed[1411],seed[729],seed[3295],seed[3804],seed[2755],seed[3758],seed[345],seed[1092],seed[2115],seed[38],seed[3788],seed[2780],seed[615],seed[376],seed[2335],seed[2405],seed[1595],seed[2441],seed[1422],seed[1874],seed[2536],seed[1950],seed[3187],seed[1522],seed[3701],seed[4002],seed[2297],seed[1803],seed[320],seed[1687],seed[4080],seed[167],seed[361],seed[2567],seed[2629],seed[3328],seed[87],seed[3754],seed[518],seed[1403],seed[897],seed[50],seed[469],seed[2692],seed[1881],seed[3062],seed[1724],seed[1063],seed[3147],seed[3666],seed[1421],seed[504],seed[472],seed[3538],seed[505],seed[1483],seed[2891],seed[284],seed[4029],seed[195],seed[2974],seed[3263],seed[4077],seed[1440],seed[3968],seed[762],seed[2577],seed[2608],seed[3422],seed[2797],seed[57],seed[3856],seed[53],seed[3104],seed[756],seed[468],seed[2654],seed[2522],seed[1868],seed[3469],seed[279],seed[1223],seed[3894],seed[3774],seed[278],seed[1733],seed[459],seed[560],seed[379],seed[303],seed[2480],seed[2049],seed[3386],seed[2526],seed[3801],seed[3324],seed[3419],seed[1509],seed[2564],seed[1710],seed[631],seed[2386],seed[3813],seed[3559],seed[1257],seed[3565],seed[981],seed[1457],seed[817],seed[1301],seed[1132],seed[2002],seed[3343],seed[3159],seed[1995],seed[3488],seed[859],seed[2326],seed[1618],seed[1906],seed[1359],seed[1073],seed[1443],seed[373],seed[3911],seed[3983],seed[3473],seed[1495],seed[3999],seed[2006],seed[719],seed[3859],seed[325],seed[686],seed[1716],seed[2980],seed[714],seed[1084],seed[3264],seed[3352],seed[3920],seed[425],seed[235],seed[3748],seed[3716],seed[3004],seed[3305],seed[1600],seed[1485],seed[1241],seed[1978],seed[354],seed[559],seed[1972],seed[3050],seed[280],seed[1946],seed[3568],seed[751],seed[3790],seed[1012],seed[1988],seed[1860],seed[887],seed[2309],seed[349],seed[1944],seed[481],seed[3331],seed[3183],seed[1127],seed[3327],seed[1051],seed[3358],seed[1765],seed[1222],seed[2303],seed[1956],seed[2788],seed[1294],seed[3811],seed[728],seed[713],seed[2734],seed[939],seed[2594],seed[445],seed[705],seed[2603],seed[3762],seed[1192],seed[498],seed[3923],seed[910],seed[944],seed[10],seed[2599],seed[471],seed[1214],seed[1052],seed[2321],seed[3065],seed[977],seed[2631],seed[989],seed[1243],seed[2410],seed[2378],seed[3550],seed[2904],seed[2293],seed[1939],seed[2794],seed[1774],seed[1409],seed[281],seed[45],seed[1809],seed[2440],seed[663],seed[3532],seed[26],seed[1410],seed[894],seed[2957],seed[1478],seed[246],seed[1463],seed[2659],seed[3945],seed[1932],seed[1702],seed[2394],seed[2031],seed[904],seed[2357],seed[2077],seed[517],seed[1402],seed[3092],seed[3600],seed[3592],seed[241],seed[1374],seed[3392],seed[1689],seed[2497],seed[2197],seed[125],seed[3980],seed[2459],seed[405],seed[1959],seed[3868],seed[3006],seed[1417],seed[1632],seed[3761],seed[2381],seed[119],seed[1905],seed[388],seed[1549],seed[122],seed[1908],seed[309],seed[2337],seed[3049],seed[1725],seed[2512],seed[3020],seed[785],seed[406],seed[610],seed[537],seed[2464],seed[3306],seed[750],seed[2126],seed[2073],seed[2258],seed[3749],seed[2889],seed[3776],seed[699],seed[2754],seed[886],seed[1130],seed[2703],seed[301],seed[56],seed[174],seed[2856],seed[37],seed[2655],seed[1255],seed[1165],seed[1302],seed[2924],seed[17],seed[2746],seed[1379],seed[1900],seed[172],seed[1866],seed[434],seed[2552],seed[2485],seed[942],seed[3582],seed[1796],seed[644],seed[2284],seed[1547],seed[973],seed[2361],seed[914],seed[742],seed[131],seed[1569],seed[3099],seed[3955],seed[1178],seed[2105],seed[2510],seed[3432],seed[621],seed[2963],seed[854],seed[1518],seed[3090],seed[3756],seed[2084],seed[2032],seed[2778],seed[232],seed[3470],seed[2622],seed[1247],seed[1129],seed[3985],seed[446],seed[3970],seed[2684],seed[820],seed[3074],seed[2779],seed[3026],seed[834],seed[2408],seed[3881],seed[2358],seed[2146],seed[1033],seed[1098],seed[24],seed[1358],seed[1365],seed[576],seed[3862],seed[2059],seed[2202],seed[2030],seed[264],seed[3739],seed[2286],seed[1631],seed[2467],seed[2819],seed[3408],seed[1591],seed[2866],seed[3782],seed[2717],seed[2356],seed[2667],seed[3512],seed[658],seed[1471],seed[3892],seed[1388],seed[1008],seed[3083],seed[4001],seed[1321],seed[3322],seed[1057],seed[1311],seed[3082],seed[3908],seed[441],seed[3043],seed[1590],seed[3040],seed[2620],seed[3864],seed[3848],seed[477],seed[1880],seed[2353],seed[1987],seed[3665],seed[930],seed[1544],seed[1465],seed[3721],seed[664],seed[247],seed[3037],seed[3845],seed[110],seed[1315],seed[3188],seed[4090],seed[83],seed[128],seed[3723],seed[860],seed[3553],seed[66],seed[557],seed[838],seed[563],seed[3109],seed[1164],seed[2498],seed[3566],seed[3335],seed[3141],seed[1851],seed[1775],seed[409],seed[3198],seed[1914],seed[2219],seed[99],seed[1248],seed[488],seed[1751],seed[1316],seed[3373],seed[532],seed[287],seed[578],seed[1496],seed[3610],seed[2148],seed[1034],seed[265],seed[3866],seed[754],seed[898],seed[2587],seed[2149],seed[3735],seed[2513],seed[3024],seed[2796],seed[1447],seed[29],seed[1286],seed[2461],seed[1917],seed[3885],seed[1427],seed[1657],seed[3533],seed[1021],seed[1264],seed[3240],seed[2199],seed[3991],seed[1455],seed[1579],seed[451],seed[2504],seed[20],seed[2768],seed[1611],seed[156],seed[2132],seed[3265],seed[3226],seed[2832],seed[3303],seed[1307],seed[3310],seed[1991],seed[3193],seed[3094],seed[1267],seed[3140],seed[1329],seed[3564],seed[3114],seed[2117],seed[3562],seed[2183],seed[873],seed[1965],seed[1607],seed[2785],seed[259],seed[2065],seed[799],seed[2244],seed[1167],seed[62],seed[1690],seed[3919],seed[1971],seed[3658],seed[2984],seed[948],seed[765],seed[3354],seed[2726],seed[643],seed[2041],seed[1501],seed[2990],seed[1259],seed[3677],seed[2831],seed[191],seed[4091],seed[1090],seed[1545],seed[760],seed[701],seed[2211],seed[4086],seed[42],seed[2813],seed[2596],seed[2666],seed[3942],seed[1011],seed[825],seed[923],seed[2938],seed[3871],seed[2660],seed[1378],seed[462],seed[3551],seed[1933],seed[3249],seed[1249],seed[4041],seed[801],seed[779],seed[4078],seed[47],seed[2881],seed[1295],seed[3606],seed[1135],seed[3046],seed[3100],seed[199],seed[826],seed[1854],seed[2157],seed[2822],seed[1674],seed[294],seed[3172],seed[1548],seed[3047],seed[2875],seed[2078],seed[2589],seed[3819],seed[1628],seed[2442],seed[3715],seed[2068],seed[1076],seed[2652],seed[386],seed[2960],seed[3587],seed[63],seed[2772],seed[41],seed[2676],seed[450],seed[1490],seed[109],seed[306],seed[2252],seed[691],seed[3405],seed[366],seed[534],seed[1145],seed[3662],seed[3398],seed[1969],seed[2551],seed[1675],seed[1508],seed[2245],seed[1213],seed[256],seed[1094],seed[608],seed[3858],seed[3279],seed[368],seed[2989],seed[3717],seed[1512],seed[1562],seed[3725],seed[2952],seed[1152],seed[2045],seed[815],seed[2349],seed[2167],seed[938],seed[3337],seed[3447],seed[3729],seed[960],seed[302],seed[190],seed[2827],seed[1584],seed[1640],seed[702],seed[203],seed[726],seed[2354],seed[3732],seed[793],seed[2396],seed[3524],seed[879],seed[795],seed[2886],seed[2109],seed[3444],seed[3572],seed[851],seed[707],seed[48],seed[3602],seed[229],seed[3318],seed[3613],seed[2277],seed[2592],seed[2259],seed[1003],seed[3428],seed[3989],seed[2131],seed[1819],seed[347],seed[2083],seed[3841],seed[2023],seed[1361],seed[2830],seed[571],seed[3687],seed[2092],seed[911],seed[221],seed[1536],seed[3575],seed[463],seed[3403],seed[2330],seed[3150],seed[1790],seed[1350],seed[496],seed[2],seed[3072],seed[4028],seed[722],seed[455],seed[1139],seed[1177],seed[3771],seed[3796],seed[3863],seed[1131],seed[2384],seed[2686],seed[2748],seed[217],seed[1760],seed[1059],seed[2409],seed[1029],seed[1753],seed[2093],seed[1990],seed[3088],seed[1338],seed[890],seed[2393],seed[3805],seed[2067],seed[314],seed[3259],seed[556],seed[3926],seed[3620],seed[3767],seed[2194],seed[1191],seed[1945],seed[3077],seed[3590],seed[568],seed[1525],seed[3946],seed[1170],seed[433],seed[142],seed[3630],seed[1438],seed[3569],seed[2176],seed[1231],seed[4055],seed[1610],seed[3807],seed[2407],seed[2472],seed[1567],seed[3786],seed[1656],seed[524],seed[551],seed[15],seed[3397],seed[1458],seed[1817],seed[408],seed[151],seed[414],seed[3329],seed[2075],seed[263],seed[2417],seed[2269],seed[3938],seed[3728],seed[2085],seed[3873],seed[3054],seed[393],seed[584],seed[3842],seed[2925],seed[3144],seed[1185],seed[3194],seed[3675],seed[2809],seed[28],seed[3297],seed[2168],seed[1718],seed[1493],seed[255],seed[995],seed[2908],seed[602],seed[2360],seed[1048],seed[2020],seed[2029],seed[2742],seed[3791],seed[2968],seed[4022],seed[979],seed[2207],seed[639],seed[1309],seed[1186],seed[1091],seed[2366],seed[1107],seed[118],seed[1028],seed[1621],seed[1001],seed[3402],seed[2022],seed[3173],seed[1744],seed[149],seed[2420],seed[1531],seed[159],seed[3168],seed[4069],seed[1182],seed[2229],seed[1682],seed[2400],seed[2475],seed[2155],seed[1892],seed[1303],seed[2364],seed[137],seed[2907],seed[2350],seed[3401],seed[1712],seed[508],seed[3434],seed[2003],seed[102],seed[359],seed[1000],seed[1190],seed[4013],seed[3288],seed[1752],seed[3940],seed[3657],seed[2451],seed[2541],seed[2833],seed[866],seed[2661],seed[1380],seed[3850],seed[1520],seed[4047],seed[478],seed[2545],seed[2088],seed[1616],seed[943],seed[842],seed[1613],seed[968],seed[2962],seed[3986],seed[2341],seed[1366],seed[3686],seed[283],seed[5],seed[2557],seed[2910],seed[1873],seed[3482],seed[3356],seed[1916],seed[3361],seed[2005],seed[2853],seed[227],seed[1810],seed[1570],seed[2205],seed[3124],seed[3959],seed[1273],seed[3884],seed[3051],seed[2715],seed[3022],seed[2195],seed[2142],seed[525],seed[3847],seed[3376],seed[470],seed[976],seed[1808],seed[3583],seed[2431],seed[2130],seed[1553],seed[2502],seed[411],seed[2678],seed[635],seed[603],seed[1814],seed[1878],seed[3627],seed[2274],seed[2438],seed[3477],seed[1435],seed[3531],seed[1327],seed[2773],seed[64],seed[3253],seed[2333],seed[1699],seed[3233],seed[3336],seed[741],seed[1849],seed[3816],seed[1523],seed[2285],seed[3446],seed[1439],seed[58],seed[1749],seed[3417],seed[1842],seed[3547],seed[3918],seed[3181],seed[1957],seed[1256],seed[484],seed[2385],seed[3759],seed[3388],seed[1179],seed[2818],seed[4021],seed[1862],seed[3586],seed[2816],seed[3423],seed[3084],seed[240],seed[1449],seed[3780],seed[213],seed[3646],seed[493],seed[2931],seed[3034],seed[464],seed[1821],seed[2267],seed[86],seed[630],seed[3400],seed[2540],seed[1331],seed[3413],seed[298],seed[296],seed[2680],seed[945],seed[3890],seed[864],seed[1277],seed[267],seed[3746],seed[3680],seed[1961],seed[2930],seed[2912],seed[2793],seed[1089],seed[3087],seed[2340],seed[2403],seed[2812],seed[2013],seed[126],seed[3979],seed[1300],seed[1346],seed[1150],seed[2255],seed[1585],seed[1187],seed[3653],seed[1464],seed[1634],seed[1037],seed[2642],seed[1505],seed[899],seed[2479],seed[1499],seed[3963],seed[2111],seed[3793],seed[339],seed[1895],seed[1183],seed[882],seed[3229],seed[1103],seed[3317],seed[2991],seed[2578],seed[1620],seed[3439],seed[1401],seed[3997],seed[2842],seed[4087],seed[3710],seed[16],seed[30],seed[3255],seed[922],seed[2489],seed[237],seed[790],seed[3891],seed[4026],seed[3299],seed[1289],seed[2374],seed[439],seed[2008],seed[852],seed[1676],seed[1383],seed[2581],seed[395],seed[1535],seed[2864],seed[4059],seed[304],seed[132],seed[1460],seed[3992],seed[313],seed[1831],seed[1587],seed[3849],seed[100],seed[4081],seed[687],seed[2492],seed[1811],seed[3511],seed[1369],seed[3014],seed[1723],seed[949],seed[2591],seed[3117],seed[44],seed[2995],seed[176],seed[1437],seed[1912],seed[2543],seed[2064],seed[419],seed[454],seed[3492],seed[1708],seed[1521],seed[1847],seed[3574],seed[2439],seed[1047],seed[3611],seed[3236],seed[2714],seed[2137],seed[2500],seed[1386],seed[428],seed[2081],seed[2346],seed[2763],seed[249],seed[260],seed[1729],seed[2369],seed[269],seed[3218],seed[582],seed[2644],seed[757],seed[3977],seed[2588],seed[2877],seed[2234],seed[3964],seed[1334],seed[1283],seed[905],seed[1915],seed[2242],seed[3817],seed[2455],seed[2736],seed[1233],seed[2936],seed[2690],seed[2488],seed[581],seed[3778],seed[1896],seed[1351],seed[348],seed[3016],seed[1859],seed[1227],seed[783],seed[3179],seed[810],seed[2272],seed[3844],seed[1020],seed[2430],seed[591],seed[613],seed[1822],seed[4093],seed[1344],seed[4044],seed[2352],seed[2021],seed[2074],seed[1189],seed[2909],seed[2294],seed[3038],seed[1577],seed[2579],seed[1111],seed[3001],seed[1042],seed[619],seed[3132],seed[650],seed[2169],seed[3041],seed[1099],seed[2201],seed[2313],seed[2494],seed[78],seed[3537],seed[2230],seed[3763],seed[818],seed[2981],seed[3585],seed[926],seed[4037],seed[97],seed[660],seed[92],seed[855],seed[401],seed[3895],seed[2870],seed[1973],seed[3852],seed[903],seed[928],seed[1080],seed[1596],seed[917],seed[2390],seed[1588],seed[3378],seed[1839],seed[494],seed[2299],seed[2628],seed[3426],seed[3390],seed[611],seed[836],seed[2977],seed[739],seed[3549],seed[2150],seed[2840],seed[1426],seed[2979],seed[2082],seed[1196],seed[3010],seed[3015],seed[3308],seed[1125],seed[3081],seed[2720],seed[2911],seed[2036],seed[3594],seed[2807],seed[2988],seed[787],seed[2215],seed[396],seed[1533],seed[3381],seed[1719],seed[2550],seed[1149],seed[2943],seed[1804],seed[372],seed[2964],seed[2921],seed[4038],seed[3523],seed[473],seed[27],seed[1756],seed[3121],seed[1335],seed[1216],seed[3563],seed[166],seed[288],seed[2711],seed[3867],seed[1172],seed[1857],seed[307],seed[2416],seed[2397],seed[2572],seed[3802],seed[402],seed[1864],seed[1260],seed[242],seed[2733],seed[3466],seed[479],seed[768],seed[3738],seed[2836],seed[1055],seed[1633],seed[2343],seed[2537],seed[3768],seed[3212],seed[2917],seed[627],seed[2610],seed[3205],seed[188],seed[2586],seed[920],seed[1560],seed[3752],seed[870],seed[1328],seed[1899],seed[1843],seed[1066],seed[858],seed[1664],seed[290],seed[1475],seed[173],seed[593],seed[1700],seed[2329],seed[1479],seed[2902],seed[2476],seed[3190],seed[1370],seed[720],seed[70],seed[3810],seed[3984],seed[1313],seed[3903],seed[3684],seed[1832],seed[2138],seed[992],seed[1732],seed[2331],seed[2424],seed[3522],seed[3461],seed[1392],seed[1825],seed[14],seed[3837],seed[1647],seed[2719],seed[3973],seed[878],seed[1109],seed[3133],seed[2009],seed[1638],seed[1606],seed[3750],seed[3091],seed[4011],seed[22],seed[2217],seed[1938],seed[1156],seed[321],seed[3883],seed[274],seed[1788],seed[839],seed[500],seed[1054],seed[622],seed[3449],seed[558],seed[1979],seed[3196],seed[2198],seed[802],seed[2898],seed[2555],seed[3468],seed[2163],seed[2287],seed[2054],seed[3822],seed[380],seed[1798],seed[2783],seed[3019],seed[72],seed[2445],seed[1105],seed[913],seed[717],seed[79],seed[1472],seed[513],seed[753],seed[4073],seed[1355],seed[1764],seed[1219],seed[3334],seed[777],seed[1703],seed[3475],seed[1714],seed[2569],seed[2934],seed[3418],seed[1356],seed[2289],seed[1993],seed[1262],seed[218],seed[3452],seed[2239],seed[238],seed[2000],seed[134],seed[2829],seed[194],seed[3474],seed[1412],seed[2119],seed[2519],seed[3244],seed[3953],seed[1685],seed[387],seed[2602],seed[3399],seed[1780],seed[3902],seed[620],seed[4085],seed[1861],seed[2246],seed[3624],seed[7],seed[752],seed[3679],seed[3900],seed[3459],seed[1787],seed[1481],seed[2791],seed[1888],seed[772],seed[3456],seed[2200],seed[933],seed[3230],seed[3301],seed[3250],seed[638],seed[3650],seed[3165],seed[1252],seed[1341],seed[3185],seed[2270],seed[577],seed[75],seed[3228],seed[3321],seed[1395],seed[3266],seed[1801],seed[3048],seed[1199],seed[3239],seed[1722],seed[3577],seed[1797],seed[2658],seed[671],seed[3286],seed[2300],seed[543],seed[2276],seed[3129],seed[1433],seed[2525],seed[2982],seed[2883],seed[2177],seed[3588],seed[1741],seed[0],seed[2641],seed[711],seed[636],seed[3772],seed[1925],seed[11],seed[4084],seed[421],seed[2486],seed[1599],seed[3861],seed[3031],seed[1038],seed[936],seed[970],seed[1602],seed[1581],seed[1642],seed[1923],seed[1017],seed[2491],seed[3812],seed[954],seed[3834],seed[3023],seed[2110],seed[1070],seed[614],seed[226],seed[1235],seed[1237],seed[998],seed[3875],seed[2709],seed[272],seed[1662],seed[1418],seed[694],seed[2933],seed[3383],seed[1065],seed[3654],seed[2638],seed[1002],seed[1404],seed[3106],seed[2878],seed[2481],seed[2266],seed[3939],seed[3311],seed[91],seed[1646],seed[123],seed[3319],seed[346],seed[625],seed[1220],seed[3056],seed[552],seed[2520],seed[1608],seed[2976],seed[3741],seed[165],seed[2640],seed[2528],seed[2634],seed[849],seed[2670],seed[3170],seed[1360],seed[2745],seed[3534],seed[609],seed[2969],seed[1290],seed[334],seed[2739],seed[168],seed[1119],seed[1261],seed[4031],seed[2249],seed[3612],seed[2688],seed[3818],seed[2428],seed[1942],seed[1100],seed[32],seed[2694],seed[1128],seed[480],seed[1693],seed[1727],seed[1684],seed[606],seed[670],seed[1820],seed[2511],seed[1171],seed[3030],seed[3874],seed[974],seed[1879],seed[586],seed[214],seed[3663],seed[1434],seed[2241],seed[1476],seed[1603],seed[353],seed[197],seed[1030],seed[3672],seed[2070],seed[343],seed[3690],seed[776],seed[1342],seed[2553],seed[3860],seed[2433],seed[3993],seed[587],seed[3478],seed[3357],seed[3651],seed[983],seed[3674],seed[940],seed[3118],seed[2291],seed[1678],seed[1343],seed[3623],seed[3581],seed[385],seed[901],seed[1557],seed[1853],seed[3536],seed[3541],seed[835],seed[963],seed[966],seed[1967],seed[812],seed[3269],seed[3634],seed[3580],seed[2371],seed[3184],seed[1598],seed[3167],seed[1511],seed[2539],seed[328],seed[3192],seed[3070],seed[3508],seed[1755],seed[2611],seed[4018],seed[2388],seed[773],seed[3377],seed[3227],seed[3348],seed[3201],seed[2687],seed[3427],seed[1113],seed[3130],seed[642],seed[2037],seed[2697],seed[3896],seed[2404],seed[895],seed[1568],seed[828],seed[317],seed[607],seed[1738],seed[397],seed[185],seed[2112],seed[3374],seed[1743],seed[330],seed[3008],seed[121],seed[3120],seed[791],seed[1492],seed[146],seed[1391],seed[1966],seed[4070],seed[1203],seed[1924],seed[2209],seed[2190],seed[152],seed[1240],seed[427],seed[497],seed[2173],seed[2418],seed[4075],seed[1445],seed[1234],seed[1834],seed[3988],seed[2087],seed[490],seed[1450],seed[4074],seed[1566],seed[3142],seed[1502],seed[1828],seed[148],seed[3839],seed[600],seed[3929],seed[962],seed[659],seed[1477],seed[1175],seed[2204],seed[270],seed[2237],seed[323],seed[3096],seed[2164],seed[646],seed[3671],seed[257],seed[1707],seed[975],seed[626],seed[1332],seed[3174],seed[2873],seed[2800],seed[426],seed[2338],seed[1800],seed[2421],seed[2236],seed[2063],seed[1058],seed[3698],seed[3209],seed[544],seed[461],seed[2834],seed[1202],seed[2452],seed[3597],seed[2328],seed[3713],seed[1265],seed[3448],seed[326],seed[2129],seed[475],seed[3075],seed[655],seed[2517],seed[1486],seed[3670],seed[3846],seed[1555],seed[4043],seed[437],seed[483],seed[3972],seed[1032],seed[2534],seed[2787],seed[3497],seed[1056],seed[3708],seed[4009],seed[3119],seed[3290],seed[845],seed[2225],seed[925],seed[3969],seed[252],seed[3640],seed[2767],seed[3578],seed[3143],seed[3649],seed[889],seed[755],seed[3262],seed[2345],seed[589],seed[3287],seed[1806],seed[1372],seed[3783],seed[3510],seed[209],seed[186],seed[1982],seed[1921],seed[3800],seed[3952],seed[2166],seed[273],seed[3136],seed[3216],seed[3450],seed[1763],seed[2508],seed[2247],seed[2264],seed[1672],seed[1487],seed[792],seed[3806],seed[352],seed[1594],seed[2696],seed[3699],seed[703],seed[3694],seed[2228],seed[3760],seed[436],seed[1060],seed[3214],seed[1556],seed[2636],seed[892],seed[2590],seed[3298],seed[1345],seed[4034],seed[3393],seed[171],seed[258],seed[2605],seed[616],seed[95],seed[391],seed[3498],seed[3080],seed[1115],seed[4066],seed[381],seed[3916],seed[1120],seed[2626],seed[3409],seed[1044],seed[3529],seed[2771],seed[1158],seed[1193],seed[2633],seed[2103],seed[2630],seed[3221],seed[3155],seed[1726],seed[3005],seed[3],seed[1102],seed[3242],seed[2178],seed[3703],seed[1325],seed[3976],seed[3154],seed[1340],seed[2625],seed[2339],seed[999],seed[189],seed[651],seed[71],seed[245],seed[90],seed[3044],seed[2133],seed[3176],seed[1292],seed[1067],seed[3616],seed[3355],seed[204],seed[3163],seed[1903],seed[1242],seed[1552],seed[363],seed[997],seed[2033],seed[2732],seed[1166],seed[2443],seed[3573],seed[1563],seed[3887],seed[1104],seed[2826],seed[1571],seed[2531],seed[3705],seed[94],seed[1393],seed[803],seed[514],seed[2320],seed[1737],seed[2436],seed[192],seed[3455],seed[2454],seed[355],seed[3851],seed[3058],seed[1592],seed[668],seed[647],seed[2055],seed[1491],seed[18],seed[2124],seed[1936],seed[3364],seed[1735],seed[3539],seed[300],seed[1144],seed[3922],seed[35],seed[1695],seed[362],seed[2501],seed[2256],seed[1937],seed[268],seed[676],seed[1748],seed[3530],seed[1474],seed[3105],seed[3639],seed[2446],seed[1123],seed[3467],seed[1155],seed[3256],seed[181],seed[2784],seed[738],seed[2248],seed[1671],seed[61],seed[813],seed[1734],seed[725],seed[683],seed[3645],seed[2056],seed[3487],seed[2095],seed[2317],seed[769],seed[1901],seed[1885],seed[3501],seed[2915],seed[1835],seed[4012],seed[1742],seed[2001],seed[3280],seed[2414],seed[1597],seed[2507],seed[1217],seed[906],seed[1406],seed[3182],seed[950],seed[1992],seed[3625],seed[3779],seed[3442],seed[3098],seed[3787],seed[1333],seed[782],seed[2387],seed[3935],seed[681],seed[2691],seed[3283],seed[3384],seed[2559],seed[1306],seed[1271],seed[2262],seed[443],seed[2187],seed[978],seed[2774],seed[2156],seed[3210],seed[3292],seed[2724],seed[3372],seed[654],seed[3349],seed[3681],seed[1337],seed[1653],seed[1413],seed[1253],seed[3309],seed[3103],seed[1462],seed[360],seed[116],seed[4],seed[3350],seed[2897],seed[2945],seed[2524],seed[1444],seed[526],seed[377],seed[503],seed[2882],seed[1244],seed[2677],seed[3367],seed[3435],seed[2435],seed[458],seed[667],seed[2325],seed[1124],seed[1210],seed[1526],seed[2972],seed[2468],seed[447],seed[2399],seed[2530],seed[3949],seed[2254],seed[1362],seed[2913],seed[3833],seed[2509],seed[2682],seed[327],seed[1229],seed[1540],seed[1539],seed[2458],seed[2208],seed[145],seed[2144],seed[356],seed[2604],seed[3491],seed[1218],seed[2025],seed[1534],seed[3353],seed[2425],seed[179],seed[383],seed[432],seed[2226],seed[3460],seed[2066],seed[3248],seed[3064],seed[1024],seed[3961],seed[3425],seed[3730],seed[1681],seed[2741],seed[2942],seed[692],seed[3500],seed[2465],seed[3344],seed[1953],seed[1083],seed[3463],seed[3893],seed[1644],seed[2948],seed[2810],seed[3669],seed[2985],seed[3203],seed[3029],seed[1405],seed[2858],seed[3486],seed[1200],seed[1468],seed[3514],seed[931],seed[2849],seed[766],seed[3965],seed[535],seed[3441],seed[412],seed[2848],seed[3584],seed[3177],seed[474],seed[3808],seed[33],seed[3134],seed[876],seed[133],seed[3371],seed[3794],seed[1280],seed[3282],seed[3489],seed[3270],seed[2304],seed[2456],seed[1758],seed[3656],seed[2868],seed[1087]}; 
//        seed3 <= {seed[1918],seed[524],seed[3736],seed[2813],seed[199],seed[1877],seed[299],seed[1459],seed[3365],seed[1019],seed[550],seed[1652],seed[1815],seed[3082],seed[2685],seed[1261],seed[2778],seed[269],seed[1253],seed[710],seed[1408],seed[506],seed[3304],seed[3540],seed[4075],seed[3862],seed[3824],seed[2929],seed[3322],seed[1474],seed[1719],seed[1929],seed[940],seed[1973],seed[3816],seed[2149],seed[725],seed[3755],seed[2172],seed[572],seed[408],seed[1939],seed[607],seed[1956],seed[2419],seed[1892],seed[2129],seed[2101],seed[1917],seed[3835],seed[3552],seed[1433],seed[1429],seed[1205],seed[1716],seed[2193],seed[2287],seed[3668],seed[4050],seed[3993],seed[2092],seed[1188],seed[544],seed[585],seed[2808],seed[3687],seed[1507],seed[641],seed[1916],seed[2469],seed[2726],seed[3726],seed[1197],seed[3228],seed[870],seed[3520],seed[1931],seed[3600],seed[2661],seed[2875],seed[2632],seed[2576],seed[3371],seed[1386],seed[3264],seed[63],seed[1338],seed[2128],seed[1496],seed[1828],seed[2691],seed[2373],seed[221],seed[952],seed[4048],seed[4044],seed[289],seed[3339],seed[1935],seed[1388],seed[2806],seed[189],seed[875],seed[4014],seed[447],seed[336],seed[1802],seed[2209],seed[384],seed[1218],seed[2985],seed[3451],seed[1641],seed[169],seed[1219],seed[1048],seed[1660],seed[713],seed[2820],seed[201],seed[3970],seed[1453],seed[1961],seed[1899],seed[1689],seed[3751],seed[2647],seed[900],seed[2842],seed[3455],seed[3899],seed[3914],seed[3605],seed[1572],seed[1708],seed[1469],seed[172],seed[3599],seed[37],seed[2038],seed[1791],seed[1749],seed[87],seed[1411],seed[2925],seed[1810],seed[2178],seed[534],seed[559],seed[1413],seed[2219],seed[1770],seed[797],seed[1982],seed[1706],seed[1595],seed[1705],seed[3399],seed[3139],seed[520],seed[3284],seed[1694],seed[3386],seed[565],seed[2447],seed[1299],seed[2829],seed[3793],seed[3700],seed[2918],seed[946],seed[3472],seed[1430],seed[2708],seed[3784],seed[263],seed[1883],seed[3693],seed[2672],seed[3996],seed[1552],seed[2170],seed[2237],seed[3646],seed[1966],seed[3643],seed[795],seed[1486],seed[1500],seed[467],seed[344],seed[1070],seed[3978],seed[3189],seed[3468],seed[2010],seed[3044],seed[2114],seed[3525],seed[1331],seed[3799],seed[1896],seed[3030],seed[4000],seed[3895],seed[3249],seed[883],seed[2700],seed[3613],seed[101],seed[1067],seed[3321],seed[874],seed[910],seed[2338],seed[2014],seed[3579],seed[1290],seed[3880],seed[906],seed[4043],seed[3967],seed[1281],seed[3834],seed[3923],seed[3063],seed[951],seed[2159],seed[1396],seed[1133],seed[329],seed[2322],seed[2750],seed[3195],seed[3889],seed[461],seed[3596],seed[2906],seed[3194],seed[1954],seed[3663],seed[3572],seed[1034],seed[1189],seed[2874],seed[3220],seed[53],seed[3795],seed[3533],seed[2481],seed[1844],seed[3404],seed[1318],seed[876],seed[3725],seed[639],seed[3919],seed[1087],seed[1555],seed[3803],seed[3577],seed[688],seed[2033],seed[3670],seed[2723],seed[2527],seed[786],seed[3746],seed[3181],seed[2085],seed[827],seed[2274],seed[1225],seed[4045],seed[252],seed[848],seed[1995],seed[2939],seed[94],seed[2834],seed[2735],seed[3580],seed[707],seed[1293],seed[3872],seed[2069],seed[2586],seed[1107],seed[3252],seed[1126],seed[3944],seed[2956],seed[208],seed[4025],seed[3973],seed[2095],seed[1049],seed[370],seed[3820],seed[3684],seed[1646],seed[2553],seed[2658],seed[122],seed[2137],seed[110],seed[148],seed[250],seed[3230],seed[2998],seed[1680],seed[1728],seed[3639],seed[1406],seed[1339],seed[3283],seed[3175],seed[1403],seed[4076],seed[1276],seed[2291],seed[2724],seed[987],seed[790],seed[1981],seed[484],seed[308],seed[1970],seed[2690],seed[115],seed[2627],seed[3591],seed[950],seed[2961],seed[989],seed[1251],seed[3859],seed[1380],seed[3361],seed[3214],seed[2802],seed[3825],seed[3818],seed[2540],seed[1834],seed[3086],seed[3901],seed[594],seed[1351],seed[3109],seed[2649],seed[1059],seed[1332],seed[2432],seed[4091],seed[2221],seed[1540],seed[497],seed[43],seed[3417],seed[1950],seed[2043],seed[3062],seed[420],seed[1495],seed[567],seed[712],seed[2631],seed[1946],seed[1988],seed[2940],seed[1588],seed[3033],seed[1300],seed[752],seed[3936],seed[1013],seed[316],seed[1710],seed[1359],seed[369],seed[3647],seed[2602],seed[1852],seed[1887],seed[2339],seed[2155],seed[3683],seed[3458],seed[1608],seed[3958],seed[4090],seed[719],seed[241],seed[501],seed[1817],seed[3087],seed[185],seed[2119],seed[3509],seed[2],seed[652],seed[3383],seed[2941],seed[2667],seed[2390],seed[2046],seed[1944],seed[2548],seed[3966],seed[3989],seed[2427],seed[334],seed[637],seed[1444],seed[3065],seed[2888],seed[3446],seed[967],seed[2426],seed[3499],seed[3794],seed[2465],seed[3199],seed[574],seed[805],seed[2721],seed[311],seed[895],seed[464],seed[2276],seed[3396],seed[616],seed[3720],seed[3701],seed[538],seed[3301],seed[3166],seed[3257],seed[3131],seed[1236],seed[3573],seed[1229],seed[1230],seed[291],seed[2972],seed[2747],seed[292],seed[1745],seed[3001],seed[2135],seed[4006],seed[1357],seed[1704],seed[3436],seed[1523],seed[728],seed[1957],seed[1363],seed[1120],seed[1860],seed[4060],seed[1836],seed[1135],seed[1978],seed[1057],seed[621],seed[2551],seed[2230],seed[2899],seed[166],seed[1132],seed[936],seed[2120],seed[4047],seed[3717],seed[2962],seed[1266],seed[4092],seed[434],seed[1687],seed[3928],seed[2526],seed[3084],seed[379],seed[1161],seed[153],seed[4023],seed[774],seed[1930],seed[1894],seed[3187],seed[824],seed[1167],seed[3739],seed[1345],seed[2652],seed[3129],seed[1808],seed[74],seed[1594],seed[2454],seed[1385],seed[2885],seed[3539],seed[2964],seed[3753],seed[3363],seed[999],seed[1115],seed[38],seed[3459],seed[566],seed[2588],seed[2388],seed[1675],seed[3992],seed[1833],seed[1228],seed[1162],seed[2883],seed[1454],seed[2959],seed[1378],seed[3542],seed[3984],seed[1438],seed[2694],seed[318],seed[2025],seed[2444],seed[1280],seed[401],seed[3735],seed[613],seed[3756],seed[3217],seed[2760],seed[1233],seed[1481],seed[664],seed[2289],seed[3903],seed[2688],seed[3118],seed[3096],seed[3508],seed[1574],seed[2541],seed[1211],seed[1042],seed[2977],seed[3790],seed[3535],seed[481],seed[4008],seed[3526],seed[894],seed[3348],seed[1150],seed[3607],seed[1907],seed[1798],seed[2657],seed[3057],seed[88],seed[2697],seed[2379],seed[846],seed[1461],seed[954],seed[1544],seed[1451],seed[322],seed[355],seed[3406],seed[61],seed[210],seed[3122],seed[246],seed[2232],seed[2845],seed[2366],seed[2107],seed[3275],seed[541],seed[1110],seed[3527],seed[1457],seed[599],seed[3940],seed[3211],seed[701],seed[1392],seed[3886],seed[2909],seed[368],seed[3904],seed[2130],seed[182],seed[643],seed[2668],seed[3776],seed[2116],seed[1854],seed[96],seed[1789],seed[2403],seed[662],seed[1005],seed[2325],seed[400],seed[422],seed[2318],seed[1144],seed[1835],seed[2425],seed[3051],seed[2570],seed[2686],seed[3185],seed[3948],seed[3715],seed[3203],seed[2531],seed[1482],seed[1171],seed[86],seed[1399],seed[347],seed[124],seed[2800],seed[1725],seed[610],seed[3495],seed[290],seed[2635],seed[360],seed[2392],seed[78],seed[3375],seed[403],seed[2236],seed[3298],seed[4069],seed[2568],seed[2642],seed[1605],seed[3208],seed[668],seed[959],seed[2436],seed[3402],seed[186],seed[2995],seed[2293],seed[2294],seed[684],seed[1627],seed[3467],seed[2645],seed[3937],seed[2249],seed[321],seed[1764],seed[3150],seed[2393],seed[986],seed[1170],seed[2204],seed[1124],seed[3713],seed[3961],seed[1222],seed[3877],seed[2771],seed[676],seed[3870],seed[1422],seed[1562],seed[2165],seed[1784],seed[1800],seed[2943],seed[1296],seed[2422],seed[1409],seed[1452],seed[980],seed[1591],seed[1759],seed[861],seed[976],seed[2220],seed[33],seed[551],seed[1510],seed[1941],seed[2613],seed[3170],seed[146],seed[3100],seed[2559],seed[3123],seed[2766],seed[1282],seed[2917],seed[3390],seed[1576],seed[1185],seed[3113],seed[3716],seed[242],seed[2870],seed[3570],seed[2539],seed[4061],seed[3832],seed[837],seed[3661],seed[3916],seed[77],seed[1558],seed[305],seed[3077],seed[1116],seed[3318],seed[2983],seed[1794],seed[2757],seed[530],seed[3069],seed[836],seed[82],seed[2718],seed[1658],seed[2256],seed[111],seed[294],seed[1095],seed[2493],seed[781],seed[2184],seed[1928],seed[3838],seed[3445],seed[132],seed[812],seed[228],seed[1766],seed[921],seed[2597],seed[1182],seed[759],seed[2081],seed[964],seed[2630],seed[3733],seed[2612],seed[720],seed[1414],seed[2516],seed[3],seed[1682],seed[2368],seed[2039],seed[3632],seed[508],seed[2653],seed[2810],seed[1543],seed[2618],seed[3091],seed[2121],seed[922],seed[1448],seed[19],seed[2138],seed[1865],seed[239],seed[1200],seed[1043],seed[2755],seed[313],seed[2185],seed[1033],seed[691],seed[1686],seed[2409],seed[1653],seed[2126],seed[3206],seed[1440],seed[1202],seed[1746],seed[771],seed[4004],seed[2850],seed[222],seed[855],seed[3863],seed[3188],seed[2664],seed[1934],seed[3556],seed[1948],seed[636],seed[1097],seed[3202],seed[2903],seed[3602],seed[2103],seed[3688],seed[2681],seed[2737],seed[2509],seed[2495],seed[681],seed[6],seed[4066],seed[1822],seed[3681],seed[1436],seed[3637],seed[1437],seed[2946],seed[387],seed[730],seed[2206],seed[801],seed[474],seed[2327],seed[1164],seed[653],seed[2824],seed[2313],seed[3629],seed[978],seed[1714],seed[273],seed[749],seed[1733],seed[1175],seed[1547],seed[341],seed[2163],seed[348],seed[3172],seed[1991],seed[1602],seed[1137],seed[2110],seed[949],seed[808],seed[90],seed[3289],seed[2633],seed[3812],seed[340],seed[2926],seed[2024],seed[1927],seed[528],seed[3169],seed[4080],seed[804],seed[984],seed[729],seed[1141],seed[3448],seed[2317],seed[3505],seed[1569],seed[13],seed[1294],seed[825],seed[1659],seed[1855],seed[3900],seed[3317],seed[3089],seed[2817],seed[3822],seed[2836],seed[1045],seed[69],seed[3503],seed[3939],seed[3486],seed[1925],seed[2467],seed[1681],seed[1509],seed[1308],seed[2355],seed[452],seed[2462],seed[939],seed[1484],seed[3890],seed[1631],seed[3878],seed[767],seed[1751],seed[2345],seed[2933],seed[857],seed[934],seed[1153],seed[2947],seed[919],seed[410],seed[3130],seed[1151],seed[1667],seed[2975],seed[3652],seed[397],seed[31],seed[2458],seed[207],seed[3792],seed[3360],seed[3142],seed[3098],seed[3487],seed[2648],seed[3039],seed[1581],seed[438],seed[1499],seed[3453],seed[2329],seed[1888],seed[2854],seed[1169],seed[658],seed[1012],seed[439],seed[1367],seed[615],seed[2756],seed[2186],seed[1405],seed[376],seed[1063],seed[3427],seed[3623],seed[2793],seed[2019],seed[3857],seed[256],seed[671],seed[3247],seed[489],seed[892],seed[2240],seed[2616],seed[3915],seed[2871],seed[249],seed[3584],seed[3023],seed[3490],seed[1748],seed[721],seed[1753],seed[1598],seed[2394],seed[247],seed[2582],seed[3676],seed[365],seed[3034],seed[2740],seed[2535],seed[2518],seed[2448],seed[1382],seed[2063],seed[3235],seed[1297],seed[300],seed[204],seed[2260],seed[298],seed[3461],seed[114],seed[3642],seed[3828],seed[2936],seed[3551],seed[2594],seed[920],seed[1341],seed[1636],seed[2188],seed[4084],seed[1769],seed[1479],seed[3771],seed[1721],seed[4019],seed[1435],seed[1609],seed[2573],seed[2980],seed[1584],seed[1573],seed[3737],seed[4028],seed[1096],seed[3002],seed[457],seed[3036],seed[1007],seed[3485],seed[3645],seed[42],seed[2158],seed[3013],seed[3773],seed[1289],seed[811],seed[692],seed[58],seed[1214],seed[3968],seed[2336],seed[3450],seed[2018],seed[2272],seed[2124],seed[1355],seed[8],seed[822],seed[445],seed[3982],seed[319],seed[3059],seed[359],seed[1303],seed[1804],seed[2670],seed[2361],seed[3950],seed[64],seed[3601],seed[320],seed[1314],seed[1123],seed[869],seed[1023],seed[3161],seed[2791],seed[2468],seed[1513],seed[2797],seed[3778],seed[1824],seed[1203],seed[2253],seed[2769],seed[3581],seed[1768],seed[212],seed[3070],seed[1799],seed[3243],seed[193],seed[1397],seed[3180],seed[2752],seed[3549],seed[1945],seed[1638],seed[871],seed[2510],seed[682],seed[2026],seed[3764],seed[2442],seed[3927],seed[898],seed[2433],seed[120],seed[2315],seed[1893],seed[3798],seed[2604],seed[3564],seed[4052],seed[1348],seed[3852],seed[2037],seed[3336],seed[1320],seed[1747],seed[1587],seed[849],seed[1718],seed[2877],seed[1691],seed[3014],seed[3842],seed[1585],seed[3456],seed[192],seed[555],seed[753],seed[765],seed[744],seed[460],seed[2146],seed[1617],seed[638],seed[624],seed[2900],seed[2279],seed[3567],seed[34],seed[3072],seed[1736],seed[1535],seed[2528],seed[3775],seed[3053],seed[1254],seed[2584],seed[1343],seed[1017],seed[2581],seed[3562],seed[1387],seed[2087],seed[2572],seed[349],seed[473],seed[1467],seed[1616],seed[665],seed[2734],seed[4071],seed[3484],seed[151],seed[1996],seed[3644],seed[1078],seed[659],seed[2957],seed[3806],seed[2380],seed[202],seed[2713],seed[3494],seed[2567],seed[93],seed[686],seed[2628],seed[3514],seed[3251],seed[1058],seed[1897],seed[179],seed[2153],seed[2781],seed[2286],seed[3530],seed[740],seed[1779],seed[2994],seed[3752],seed[4081],seed[2898],seed[3449],seed[1027],seed[2076],seed[620],seed[3327],seed[1093],seed[138],seed[3424],seed[3209],seed[2514],seed[2763],seed[1047],seed[2464],seed[2320],seed[3610],seed[1538],seed[913],seed[1490],seed[2910],seed[3938],seed[3625],seed[450],seed[66],seed[3388],seed[236],seed[2984],seed[618],seed[1503],seed[449],seed[2342],seed[332],seed[220],seed[799],seed[3976],seed[2938],seed[4085],seed[4005],seed[750],seed[3179],seed[29],seed[2408],seed[3239],seed[2908],seed[1674],seed[310],seed[2386],seed[2140],seed[3529],seed[902],seed[864],seed[2682],seed[3922],seed[2494],seed[3302],seed[2415],seed[1878],seed[3557],seed[1416],seed[3658],seed[2471],seed[1163],seed[2118],seed[703],seed[1801],seed[1599],seed[3628],seed[1709],seed[1642],seed[928],seed[539],seed[1909],seed[3429],seed[1589],seed[3991],seed[2125],seed[806],seed[1391],seed[312],seed[2387],seed[1879],seed[2477],seed[134],seed[1084],seed[1707],seed[2349],seed[3924],seed[363],seed[3350],seed[3391],seed[2154],seed[492],seed[331],seed[2203],seed[1053],seed[1847],seed[1781],seed[1821],seed[2405],seed[361],seed[2347],seed[971],seed[3151],seed[2323],seed[2078],seed[260],seed[3121],seed[4030],seed[3972],seed[2701],seed[1895],seed[1076],seed[1298],seed[4059],seed[882],seed[118],seed[1842],seed[2189],seed[3691],seed[1625],seed[76],seed[3589],seed[4073],seed[1761],seed[398],seed[1172],seed[3860],seed[562],seed[431],seed[852],seed[2575],seed[746],seed[3699],seed[1943],seed[1669],seed[3017],seed[4031],seed[3430],seed[1088],seed[1178],seed[2190],seed[1863],seed[796],seed[1313],seed[1536],seed[858],seed[2466],seed[3821],seed[328],seed[2952],seed[516],seed[1183],seed[1323],seed[2622],seed[3074],seed[1922],seed[2549],seed[2222],seed[2143],seed[1592],seed[549],seed[3782],seed[2480],seed[2695],seed[3810],seed[2171],seed[3167],seed[2304],seed[3867],seed[3473],seed[788],seed[927],seed[3758],seed[2546],seed[2953],seed[3101],seed[1551],seed[3364],seed[2765],seed[1149],seed[838],seed[741],seed[28],seed[2876],seed[3474],seed[3411],seed[2057],seed[2067],seed[649],seed[734],seed[859],seed[3910],seed[2428],seed[3042],seed[1156],seed[2297],seed[3695],seed[2678],seed[1243],seed[200],seed[3397],seed[3774],seed[3696],seed[2707],seed[695],seed[1340],seed[1977],seed[2683],seed[377],seed[3447],seed[24],seed[1903],seed[3270],seed[3897],seed[209],seed[3442],seed[509],seed[2201],seed[3431],seed[2319],seed[885],seed[3544],seed[302],seed[630],seed[2932],seed[3041],seed[582],seed[3518],seed[218],seed[1241],seed[3127],seed[2866],seed[2267],seed[1419],seed[1038],seed[3560],seed[556],seed[2865],seed[2732],seed[68],seed[1514],seed[1008],seed[1328],seed[1870],seed[1002],seed[4032],seed[1985],seed[1864],seed[1624],seed[650],seed[338],seed[2555],seed[798],seed[2981],seed[2239],seed[909],seed[1545],seed[3236],seed[1434],seed[2020],seed[1035],seed[1557],seed[140],seed[3193],seed[2215],seed[961],seed[1142],seed[2282],seed[3787],seed[1426],seed[2591],seed[1011],seed[1740],seed[2410],seed[3231],seed[2411],seed[500],seed[2071],seed[3802],seed[2423],seed[1213],seed[433],seed[4013],seed[1094],seed[2292],seed[1356],seed[1867],seed[972],seed[3744],seed[850],seed[561],seed[3040],seed[3480],seed[742],seed[1190],seed[1868],seed[3233],seed[1906],seed[2086],seed[3745],seed[2229],seed[589],seed[933],seed[2132],seed[1064],seed[1085],seed[3067],seed[2809],seed[2441],seed[1654],seed[2950],seed[123],seed[1069],seed[3392],seed[1517],seed[1117],seed[3921],seed[1738],seed[1611],seed[133],seed[2619],seed[416],seed[3957],seed[1990],seed[3528],seed[1676],seed[2934],seed[2725],seed[3465],seed[1317],seed[493],seed[1677],seed[2461],seed[1284],seed[2285],seed[3641],seed[3705],seed[3075],seed[2788],seed[307],seed[3104],seed[2102],seed[14],seed[3163],seed[35],seed[2601],seed[3140],seed[3594],seed[174],seed[2484],seed[2916],seed[2307],seed[1607],seed[4036],seed[1130],seed[685],seed[3258],seed[3242],seed[119],seed[1793],seed[2060],seed[3561],seed[2712],seed[285],seed[2202],seed[2692],seed[2169],seed[3734],seed[2115],seed[3523],seed[2271],seed[4058],seed[1932],seed[581],seed[2758],seed[3708],seed[2585],seed[1335],seed[3826],seed[2547],seed[1744],seed[3489],seed[1637],seed[2344],seed[257],seed[3638],seed[2736],seed[3421],seed[1809],seed[1104],seed[2492],seed[2055],seed[3656],seed[1373],seed[588],seed[155],seed[1431],seed[1001],seed[2098],seed[3657],seed[107],seed[458],seed[2151],seed[1065],seed[57],seed[230],seed[205],seed[337],seed[40],seed[823],seed[1610],seed[1987],seed[2174],seed[1622],seed[167],seed[2210],seed[1623],seed[514],seed[1797],seed[595],seed[3016],seed[1267],seed[675],seed[648],seed[1737],seed[2655],seed[1106],seed[3918],seed[2892],seed[994],seed[1603],seed[3439],seed[2574],seed[3614],seed[3955],seed[2663],seed[975],seed[326],seed[758],seed[2283],seed[644],seed[2669],seed[766],seed[3454],seed[1796],seed[2389],seed[3300],seed[109],seed[3830],seed[814],seed[737],seed[2414],seed[2181],seed[3291],seed[1811],seed[2895],seed[718],seed[1711],seed[2812],seed[2679],seed[2557],seed[2993],seed[3340],seed[1285],seed[4093],seed[2047],seed[1235],seed[52],seed[2162],seed[3315],seed[2248],seed[2131],seed[258],seed[3931],seed[723],seed[3401],seed[3722],seed[26],seed[3709],seed[3149],seed[2006],seed[2935],seed[3056],seed[918],seed[2930],seed[633],seed[3460],seed[1920],seed[465],seed[2911],seed[2945],seed[2073],seed[5],seed[2455],seed[12],seed[1566],seed[698],seed[3960],seed[1309],seed[1006],seed[3341],seed[2357],seed[754],seed[3788],seed[2571],seed[1635],seed[2569],seed[195],seed[2815],seed[1720],seed[3706],seed[619],seed[288],seed[2218],seed[1492],seed[1952],seed[942],seed[3428],seed[1274],seed[1805],seed[270],seed[27],seed[3945],seed[444],seed[2328],seed[1021],seed[3515],seed[896],seed[309],seed[1644],seed[1795],seed[3779],seed[3232],seed[3409],seed[54],seed[1127],seed[494],seed[10],seed[571],seed[1840],seed[2879],seed[1614],seed[3005],seed[383],seed[2000],seed[352],seed[745],seed[944],seed[3225],seed[2988],seed[1307],seed[2774],seed[411],seed[1861],seed[1501],seed[904],seed[2564],seed[345],seed[2008],seed[2790],seed[1292],seed[1354],seed[2714],seed[1061],seed[583],seed[2792],seed[2265],seed[3332],seed[1962],seed[2262],seed[3178],seed[1372],seed[3124],seed[1083],seed[3303],seed[1288],seed[3833],seed[1152],seed[860],seed[275],seed[4018],seed[2651],seed[2644],seed[1633],seed[731],seed[213],seed[960],seed[2301],seed[3664],seed[1882],seed[793],seed[2872],seed[2122],seed[2108],seed[791],seed[2522],seed[3959],seed[3215],seed[2491],seed[3478],seed[3061],seed[2275],seed[59],seed[1287],seed[3675],seed[1109],seed[3543],seed[1324],seed[2023],seed[1712],seed[2029],seed[1091],seed[1407],seed[1498],seed[780],seed[2521],seed[1112],seed[2704],seed[3221],seed[1086],seed[1819],seed[3168],seed[907],seed[440],seed[1643],seed[2828],seed[611],seed[2051],seed[2263],seed[157],seed[3854],seed[1814],seed[3165],seed[1512],seed[1221],seed[3492],seed[1938],seed[2015],seed[789],seed[462],seed[3712],seed[3855],seed[1488],seed[1337],seed[569],seed[702],seed[2992],seed[0],seed[779],seed[3980],seed[164],seed[1301],seed[446],seed[1724],seed[3319],seed[2727],seed[511],seed[2839],seed[635],seed[1757],seed[603],seed[3634],seed[3942],seed[2430],seed[2331],seed[552],seed[3006],seed[1333],seed[2213],seed[2767],seed[518],seed[393],seed[3772],seed[667],seed[2924],seed[1729],seed[2278],seed[3356],seed[394],seed[1302],seed[3585],seed[196],seed[2578],seed[1255],seed[2280],seed[1304],seed[2333],seed[39],seed[3156],seed[2748],seed[997],seed[2214],seed[362],seed[844],seed[3240],seed[1311],seed[2673],seed[602],seed[2109],seed[1483],seed[1726],seed[1739],seed[3387],seed[343],seed[2965],seed[1291],seed[1604],seed[2951],seed[2354],seed[3612],seed[2141],seed[1959],seed[598],seed[3441],seed[2486],seed[1071],seed[3471],seed[2375],seed[2852],seed[1976],seed[1975],seed[1765],seed[1319],seed[3229],seed[1730],seed[1525],seed[2884],seed[3144],seed[3320],seed[3182],seed[3254],seed[628],seed[1381],seed[998],seed[2923],seed[1553],seed[1734],seed[899],seed[1515],seed[2978],seed[935],seed[760],seed[1942],seed[206],seed[925],seed[2247],seed[2782],seed[3433],seed[1018],seed[1619],seed[3029],seed[2134],seed[3164],seed[819],seed[2543],seed[265],seed[2580],seed[2050],seed[3135],seed[2905],seed[672],seed[1275],seed[18],seed[802],seed[716],seed[188],seed[223],seed[2352],seed[3674],seed[2383],seed[3907],seed[264],seed[3650],seed[2634],seed[1816],seed[3537],seed[3975],seed[3714],seed[4042],seed[1108],seed[2284],seed[1030],seed[105],seed[3218],seed[1493],seed[2300],seed[3609],seed[480],seed[1648],seed[346],seed[3197],seed[577],seed[2053],seed[3212],seed[924],seed[3060],seed[1655],seed[2893],seed[938],seed[79],seed[1081],seed[3358],seed[44],seed[2759],seed[131],seed[3586],seed[1477],seed[2840],seed[3868],seed[1803],seed[1400],seed[1999],seed[1541],seed[2048],seed[2646],seed[2034],seed[4002],seed[3250],seed[1259],seed[2517],seed[1516],seed[3416],seed[2452],seed[2127],seed[3483],seed[3626],seed[3479],seed[2823],seed[2266],seed[3248],seed[2459],seed[903],seed[1364],seed[1993],seed[3545],seed[3031],seed[2927],seed[325],seed[2536],seed[1231],seed[623],seed[415],seed[2017],seed[226],seed[3049],seed[2070],seed[219],seed[3425],seed[663],seed[2963],seed[2662],seed[564],seed[1402],seed[2420],seed[3045],seed[4034],seed[1365],seed[3174],seed[1664],seed[2506],seed[1080],seed[3521],seed[3353],seed[1131],seed[1914],seed[1068],seed[533],seed[1837],seed[1195],seed[3011],seed[884],seed[3400],seed[2890],seed[3690],seed[3136],seed[722],seed[3234],seed[3080],seed[1249],seed[2579],seed[977],seed[2715],seed[1665],seed[3437],seed[3702],seed[3742],seed[3731],seed[1898],seed[3692],seed[2948],seed[425],seed[3963],seed[979],seed[2161],seed[1165],seed[2052],seed[738],seed[1508],seed[3905],seed[600],seed[1915],seed[2478],seed[2443],seed[194],seed[1783],seed[3423],seed[1891],seed[1208],seed[259],seed[1196],seed[632],seed[1874],seed[380],seed[834],seed[2913],seed[3097],seed[2299],seed[3032],seed[2717],seed[11],seed[2421],seed[1632],seed[1775],seed[48],seed[2534],seed[1077],seed[1849],seed[3078],seed[1758],seed[3463],seed[1550],seed[553],seed[2861],seed[1082],seed[3438],seed[2321],seed[3226],seed[3892],seed[423],seed[2489],seed[2650],seed[2111],seed[2356],seed[2860],seed[2439],seed[974],seed[3493],seed[1024],seed[2722],seed[957],seed[3906],seed[3883],seed[1401],seed[3162],seed[1210],seed[2970],seed[1786],seed[941],seed[3920],seed[382],seed[3384],seed[2639],seed[1447],seed[3488],seed[626],seed[2314],seed[2805],seed[521],seed[2955],seed[1851],seed[3583],seed[1556],seed[726],seed[3640],seed[102],seed[1671],seed[2991],seed[2787],seed[931],seed[1232],seed[1806],seed[2529],seed[2498],seed[1839],seed[356],seed[2835],seed[1342],seed[476],seed[3286],seed[3055],seed[3929],seed[646],seed[95],seed[2113],seed[1845],seed[592],seed[1040],seed[841],seed[3134],seed[3048],seed[262],seed[908],seed[315],seed[2058],seed[1848],seed[593],seed[3237],seed[141],seed[1666],seed[3593],seed[3146],seed[3207],seed[631],seed[3079],seed[2391],seed[459],seed[1923],seed[3050],seed[3721],seed[3590],seed[1546],seed[3947],seed[1924],seed[498],seed[654],seed[277],seed[1717],seed[130],seed[2878],seed[968],seed[1468],seed[1240],seed[2838],seed[2590],seed[1125],seed[2777],seed[3845],seed[1394],seed[2511],seed[171],seed[2507],seed[914],seed[1020],seed[22],seed[388],seed[622],seed[49],seed[1846],seed[2479],seed[661],seed[724],seed[576],seed[266],seed[211],seed[579],seed[1361],seed[3395],seed[818],seed[2659],seed[2360],seed[2742],seed[1843],seed[1174],seed[296],seed[2770],seed[3724],seed[424],seed[2561],seed[1537],seed[1480],seed[981],seed[3550],seed[1969],seed[2921],seed[1412],seed[3502],seed[2841],seed[32],seed[2979],seed[2160],seed[1963],seed[3081],seed[3669],seed[2680],seed[3273],seed[1039],seed[1439],seed[1277],seed[2621],seed[873],seed[330],seed[1606],seed[2346],seed[3770],seed[2485],seed[3342],seed[2699],seed[4088],seed[2819],seed[178],seed[1528],seed[297],seed[3913],seed[647],seed[813],seed[4016],seed[1820],seed[2021],seed[3723],seed[3979],seed[3869],seed[170],seed[761],seed[863],seed[609],seed[2780],seed[3760],seed[1697],seed[342],seed[2863],seed[2001],seed[3804],seed[3111],seed[1158],seed[1960],seed[286],seed[1022],seed[3470],seed[700],seed[1441],seed[3413],seed[1857],seed[1889],seed[472],seed[1875],seed[2090],seed[2156],seed[679],seed[2487],seed[1521],seed[1148],seed[3815],seed[3732],seed[3635],seed[317],seed[830],seed[777],seed[504],seed[406],seed[1360],seed[739],seed[608],seed[3500],seed[1983],seed[2112],seed[2603],seed[2363],seed[512],seed[792],seed[432],seed[3837],seed[3279],seed[2552],seed[1118],seed[563],seed[3861],seed[3743],seed[85],seed[1613],seed[2512],seed[2144],seed[3685],seed[244],seed[546],seed[2438],seed[1398],seed[666],seed[1262],seed[3326],seed[2460],seed[165],seed[1621],seed[2105],seed[3337],seed[4024],seed[2503],seed[3578],seed[231],seed[1187],seed[3466],seed[2896],seed[3263],seed[3819],seed[1050],seed[333],seed[655],seed[3147],seed[3280],seed[2869],seed[1004],seed[3783],seed[4027],seed[3686],seed[3757],seed[2577],seed[2281],seed[3874],seed[2164],seed[2372],seed[3064],seed[97],seed[485],seed[2675],seed[851],seed[3844],seed[2225],seed[2592],seed[3654],seed[2401],seed[2505],seed[1559],seed[1286],seed[1979],seed[1143],seed[4077],seed[1154],seed[3606],seed[98],seed[3378],seed[3698],seed[2523],seed[1194],seed[763],seed[502],seed[1168],seed[2196],seed[1217],seed[1044],seed[2728],seed[3849],seed[3035],seed[1271],seed[1458],seed[2607],seed[36],seed[2407],seed[25],seed[2967],seed[2335],seed[2402],seed[1994],seed[3491],seed[1329],seed[1445],seed[3673],seed[3276],seed[4003],seed[1463],seed[1651],seed[350],seed[2406],seed[2440],seed[278],seed[1869],seed[2180],seed[3374],seed[727],seed[390],seed[1443],seed[1756],seed[3865],seed[3009],seed[468],seed[2605],seed[1016],seed[1427],seed[3964],seed[1327],seed[229],seed[3046],seed[2711],seed[3323],seed[1206],seed[1368],seed[3718],seed[3205],seed[1701],seed[1511],seed[2273],seed[245],seed[2986],seed[3346],seed[966],seed[2326],seed[2937],seed[1121],seed[2175],seed[2072],seed[2623],seed[3912],seed[1974],seed[683],seed[3157],seed[1936],seed[15],seed[2099],seed[2542],seed[1578],seed[191],seed[690],seed[2233],seed[2949],seed[3324],seed[956],seed[2257],seed[251],seed[2041],seed[1529],seed[1138],seed[4049],seed[2397],seed[2049],seed[893],seed[816],seed[238],seed[3971],seed[2987],seed[1315],seed[3148],seed[2556],seed[62],seed[1224],seed[2768],seed[2028],seed[2011],seed[1829],seed[1777],seed[280],seed[3385],seed[2942],seed[3648],seed[3309],seed[3563],seed[287],seed[396],seed[1727],seed[2643],seed[3373],seed[2508],seed[2194],seed[3587],seed[807],seed[443],seed[2261],seed[2089],seed[1395],seed[113],seed[3022],seed[1014],seed[3848],seed[2902],seed[3740],seed[527],seed[399],seed[3133],seed[2996],seed[2207],seed[1989],seed[3008],seed[697],seed[3839],seed[2598],seed[1580],seed[2786],seed[926],seed[2083],seed[3297],seed[2901],seed[3112],seed[142],seed[748],seed[2565],seed[568],seed[601],seed[2334],seed[2826],seed[3797],seed[4021],seed[3224],seed[1628],seed[2859],seed[2123],seed[3253],seed[3555],seed[2997],seed[1812],seed[1940],seed[421],seed[2744],seed[3840],seed[536],seed[2032],seed[3926],seed[3325],seed[2147],seed[2068],seed[696],seed[2851],seed[711],seed[3271],seed[451],seed[1871],seed[3769],seed[1257],seed[1933],seed[1362],seed[3565],seed[3592],seed[2104],seed[366],seed[3719],seed[373],seed[3780],seed[2496],seed[2638],seed[1223],seed[1683],seed[2482],seed[3186],seed[670],seed[454],seed[1560],seed[1201],seed[143],seed[2016],seed[542],seed[535],seed[2928],seed[1539],seed[958],seed[4039],seed[1593],seed[854],seed[1237],seed[1446],seed[845],seed[2044],seed[1244],seed[1853],seed[1478],seed[3536],seed[2764],seed[3697],seed[3177],seed[303],seed[3246],seed[2666],seed[2803],seed[3120],seed[3138],seed[463],seed[435],seed[3043],seed[674],seed[3891],seed[1561],seed[4035],seed[1442],seed[2502],seed[3094],seed[3210],seed[831],seed[3888],seed[2295],seed[558],seed[3941],seed[3126],seed[1542],seed[2629],seed[3310],seed[2195],seed[1565],seed[1432],seed[83],seed[116],seed[3443],seed[3379],seed[2369],seed[3152],seed[1114],seed[1866],seed[3352],seed[879],seed[2973],seed[800],seed[4087],seed[2676],seed[1713],seed[2035],seed[293],seed[3026],seed[973],seed[187],seed[364],seed[835],seed[1661],seed[3851],seed[3588],seed[3299],seed[3434],seed[4064],seed[3679],seed[2330],seed[1649],seed[3547],seed[829],seed[117],seed[2677],seed[1079],seed[890],seed[3999],seed[441],seed[3088],seed[4009],seed[2377],seed[1046],seed[2082],seed[1549],seed[3153],seed[1146],seed[2231],seed[240],seed[1754],seed[3274],seed[2912],seed[2532],seed[279],seed[1792],seed[3707],seed[1750],seed[853],seed[274],seed[2133],seed[3003],seed[1],seed[3624],seed[3879],seed[3281],seed[1404],seed[3615],seed[65],seed[2385],seed[4055],seed[327],seed[3595],seed[1173],seed[3568],seed[3766],seed[3917],seed[2378],seed[1242],seed[127],seed[1620],seed[248],seed[3076],seed[2370],seed[732],seed[768],seed[3012],seed[4020],seed[943],seed[391],seed[1346],seed[1968],seed[1100],seed[1912],seed[158],seed[2003],seed[963],seed[135],seed[3729],seed[2922],seed[306],seed[2886],seed[1807],seed[2100],seed[1533],seed[1347],seed[505],seed[108],seed[764],seed[543],seed[2814],seed[1487],seed[775],seed[982],seed[3496],seed[335],seed[1465],seed[1179],seed[3106],seed[1025],seed[3288],seed[1239],seed[150],seed[2490],seed[3930],seed[3481],seed[1475],seed[587],seed[2596],seed[499],seed[2919],seed[3951],seed[3259],seed[367],seed[3435],seed[1041],seed[3666],seed[2710],seed[2897],seed[1312],seed[2324],seed[1471],seed[235],seed[339],seed[736],seed[2862],seed[3969],seed[2264],seed[573],seed[1421],seed[1904],seed[1157],seed[3504],seed[2773],seed[1054],seed[1778],seed[3532],seed[358],seed[183],seed[2554],seed[159],seed[1826],seed[625],seed[1199],seed[1056],seed[2501],seed[2251],seed[1248],seed[2960],seed[233],seed[3285],seed[923],seed[453],seed[2277],seed[1731],seed[2030],seed[1640],seed[3018],seed[3296],seed[2907],seed[2848],seed[2858],seed[3114],seed[2625],seed[3245],seed[104],seed[983],seed[4015],seed[409],seed[173],seed[304],seed[2483],seed[3896],seed[1656],seed[1316],seed[3887],seed[3372],seed[3370],seed[3933],seed[2353],seed[1813],seed[3981],seed[3791],seed[2698],seed[2822],seed[374],seed[3864],seed[2332],seed[3498],seed[1823],seed[46],seed[1238],seed[1424],seed[3768],seed[3660],seed[2012],seed[1181],seed[1344],seed[354],seed[1696],seed[634],seed[1873],seed[1349],seed[604],seed[2614],seed[4095],seed[2772],seed[80],seed[3823],seed[3846],seed[3630],seed[1494],seed[1571],seed[2881],seed[3559],seed[3369],seed[947],seed[2079],seed[2801],seed[2013],seed[2075],seed[475],seed[2500],seed[351],seed[2362],seed[1410],seed[1155],seed[2693],seed[2418],seed[3730],seed[3636],seed[1270],seed[1204],seed[1838],seed[2191],seed[2867],seed[3137],seed[3847],seed[3811],seed[917],seed[1216],seed[699],seed[1379],seed[1715],seed[1215],seed[515],seed[1377],seed[1965],seed[3389],seed[1330],seed[1612],seed[578],seed[548],seed[3260],seed[3908],seed[3108],seed[3015],seed[1031],seed[1972],seed[517],seed[3099],seed[3415],seed[2080],seed[2600],seed[965],seed[1310],seed[3513],seed[1247],seed[2969],seed[1028],seed[2689],seed[880],seed[1191],seed[2093],seed[3125],seed[2830],seed[225],seed[3201],seed[3704],seed[3934],seed[16],seed[1634],seed[2208],seed[1752],seed[1858],seed[3665],seed[1140],seed[2847],seed[1060],seed[488],seed[2702],seed[1052],seed[856],seed[3071],seed[3198],seed[2258],seed[3512],seed[237],seed[2398],seed[785],seed[2589],seed[2416],seed[1250],seed[3393],seed[1417],seed[1072],seed[2587],seed[2544],seed[2853],seed[92],seed[1741],seed[495],seed[3954],seed[3265],seed[1489],seed[955],seed[1180],seed[1519],seed[1760],seed[1601],seed[1279],seed[522],seed[2563],seed[412],seed[2296],seed[772],seed[2197],seed[268],seed[996],seed[2417],seed[1177],seed[2891],seed[3312],seed[372],seed[2914],seed[3090],seed[2606],seed[597],seed[2234],seed[2743],seed[865],seed[1147],seed[1101],seed[3227],seed[4038],seed[3519],seed[2525],seed[203],seed[2005],seed[1524],seed[2738],seed[3255],seed[2269],seed[112],seed[378],seed[2709],seed[2413],seed[3204],seed[782],seed[3457],seed[2624],seed[3911],seed[1998],seed[1128],seed[1980],seed[4083],seed[4051],seed[2599],seed[1504],seed[1958],seed[139],seed[747],seed[3909],seed[945],seed[73],seed[3328],seed[3268],seed[1699],seed[2706],seed[2753],seed[2288],seed[2811],seed[3902],seed[353],seed[2887],seed[843],seed[629],seed[612],seed[2382],seed[371],seed[2036],seed[3349],seed[2827],seed[1009],seed[756],seed[2530],seed[1209],seed[418],seed[2303],seed[673],seed[152],seed[3667],seed[3622],seed[1567],seed[3244],seed[1672],seed[3362],seed[2227],seed[2989],seed[3680],seed[30],seed[1531],seed[2831],seed[2472],seed[3574],seed[496],seed[1911],seed[2463],seed[2641],seed[2846],seed[2312],seed[3617],seed[3813],seed[657],seed[1306],seed[3767],seed[1325],seed[2400],seed[1921],seed[2173],seed[821],seed[2562],seed[2216],seed[2719],seed[1774],seed[99],seed[3335],seed[21],seed[45],seed[3267],seed[1497],seed[2243],seed[678],seed[301],seed[2779],seed[177],seed[3266],seed[605],seed[1647],seed[2608],seed[1015],seed[2217],seed[129],seed[1971],seed[1881],seed[1722],seed[3145],seed[2894],seed[491],seed[868],seed[3477],seed[2177],seed[915],seed[3021],seed[2504],seed[3073],seed[3256],seed[1984],seed[1036],seed[163],seed[891],seed[1702],seed[106],seed[867],seed[2558],seed[161],seed[3154],seed[735],seed[1771],seed[419],seed[84],seed[1186],seed[3452],seed[3598],seed[2031],seed[1947],seed[3781],seed[3222],seed[993],seed[3403],seed[389],seed[2920],seed[2009],seed[3085],seed[1129],seed[3785],seed[136],seed[3777],seed[405],seed[3261],seed[125],seed[2311],seed[3809],seed[1010],seed[2864],seed[414],seed[803],seed[267],seed[3292],seed[4010],seed[426],seed[4001],seed[2308],seed[3190],seed[905],seed[3582],seed[2340],seed[916],seed[2615],seed[769],seed[3476],seed[1600],seed[3548],seed[1207],seed[784],seed[2179],seed[1548],seed[2749],seed[953],seed[75],seed[1520],seed[1986],seed[3807],seed[1227],seed[3377],seed[1530],seed[3619],seed[3871],seed[3678],seed[2223],seed[3893],seed[2358],seed[3338],seed[3282],seed[70],seed[3311],seed[197],seed[3765],seed[3497],seed[1832],seed[3763],seed[466],seed[1246],seed[3269],seed[3419],seed[3331],seed[3689],seed[2626],seed[4074],seed[1166],seed[3351],seed[714],seed[2091],seed[3200],seed[1755],seed[614],seed[1322],seed[3058],seed[3093],seed[198],seed[3038],seed[937],seed[1534],seed[3407],seed[833],seed[1910],seed[168],seed[2799],seed[2268],seed[4062],seed[1859],seed[1425],seed[3965],seed[2751],seed[3569],seed[2002],seed[705],seed[156],seed[3277],seed[3789],seed[2671],seed[1273],seed[2958],seed[3287],seed[1136],seed[3850],seed[470],seed[3516],seed[3994],seed[1159],seed[1780],seed[3884],seed[4086],seed[1788],seed[1418],seed[1735],seed[184],seed[3627],seed[1383],seed[2545],seed[2290],seed[2524],seed[2785],seed[540],seed[2705],seed[3501],seed[3410],seed[743],seed[1105],seed[2818],seed[751],seed[1450],seed[694],seed[385],seed[991],seed[1668],seed[3881],seed[3524],seed[2519],seed[3116],seed[1476],seed[3213],seed[2094],seed[2066],seed[1375],seed[3671],seed[2807],seed[901],seed[2637],seed[2437],seed[642],seed[3754],seed[2061],seed[2365],seed[428],seed[456],seed[4012],seed[1862],seed[3355],seed[1657],seed[1264],seed[3677],seed[911],seed[575],seed[1693],seed[2242],seed[3814],seed[1905],seed[1334],seed[3176],seed[3649],seed[1098],seed[878],seed[1937],seed[3308],seed[584],seed[455],seed[4017],seed[1506],seed[2513],seed[531],seed[1850],seed[67],seed[3946],seed[1773],seed[778],seed[2533],seed[3843],seed[3027],seed[3603],seed[2434],seed[1919],seed[3028],seed[660],seed[1670],seed[2065],seed[3511],seed[1111],seed[3531],seed[2499],seed[3128],seed[3517],seed[680],seed[1690],seed[2473],seed[2042],seed[4007],seed[284],seed[4054],seed[1700],seed[617],seed[381],seed[1522],seed[2457],seed[71],seed[704],seed[3290],seed[448],seed[2150],seed[3682],seed[2244],seed[3366],seed[1374],seed[4078],seed[2674],seed[3694],seed[733],seed[3885],seed[1762],seed[2298],seed[2849],seed[395],seed[3831],seed[930],seed[560],seed[3796],seed[1269],seed[145],seed[477],seed[2795],seed[3405],seed[3380],seed[3295],seed[794],seed[2798],seed[3998],seed[513],seed[1518],seed[877],seed[1062],seed[404],seed[1880],seed[1678],seed[3007],seed[3943],seed[3262],seed[1193],seed[3052],seed[2255],seed[1967],seed[1119],seed[3191],seed[2776],seed[554],seed[243],seed[1901],seed[783],seed[2343],seed[2364],seed[1305],seed[4046],seed[840],seed[2857],seed[3651],seed[3223],seed[606],seed[4079],seed[3988],seed[2595],seed[3749],seed[2474],seed[3949],seed[1370],seed[3054],seed[176],seed[1872],seed[3020],seed[3160],seed[2351],seed[2617],seed[645],seed[757],seed[1579],seed[2889],seed[2106],seed[2449],seed[717],seed[2609],seed[2583],seed[1688],seed[2520],seed[3805],seed[3985],seed[1350],seed[3102],seed[2904],seed[3983],seed[1134],seed[2316],seed[2739],seed[2412],seed[2445],seed[1295],seed[929],seed[651],seed[1358],seed[2976],seed[2636],seed[2399],seed[866],seed[3272],seed[1505],seed[3853],seed[2703],seed[121],seed[89],seed[1456],seed[1645],seed[3759],seed[2395],seed[1767],seed[386],seed[3728],seed[2837],seed[1890],seed[1074],seed[1663],seed[482],seed[1884],seed[2610],seed[3381],seed[689],seed[2593],seed[2730],seed[2431],seed[3738],seed[3004],seed[776],seed[3935],seed[640],seed[809],seed[557],seed[1263],seed[3105],seed[2538],seed[2429],seed[1113],seed[1145],seed[1491],seed[1420],seed[3558],seed[988],seed[656],seed[3066],seed[4053],seed[2004],seed[2816],seed[2843],seed[2982],seed[253],seed[47],seed[429],seed[2022],seed[2241],seed[1841],seed[2245],seed[1176],seed[3786],seed[3159],seed[2654],seed[2687],seed[2341],seed[4070],seed[2775],seed[3155],seed[402],seed[2833],seed[1684],seed[2376],seed[2212],seed[154],seed[2488],seed[2856],seed[708],seed[2446],seed[2371],seed[1103],seed[3898],seed[3238],seed[1787],seed[3747],seed[3829],seed[2804],seed[2096],seed[815],seed[261],seed[1732],seed[3037],seed[1390],seed[3376],seed[1856],seed[137],seed[60],seed[2784],seed[2211],seed[1597],seed[3748],seed[1055],seed[3621],seed[2224],seed[525],seed[532],seed[3987],seed[3462],seed[2270],seed[427],seed[3444],seed[479],seed[407],seed[2873],seed[3047],seed[147],seed[995],seed[669],seed[3359],seed[3095],seed[2424],seed[2306],seed[2660],seed[214],seed[2183],seed[181],seed[3952],seed[1964],seed[417],seed[2966],seed[2794],seed[828],seed[2971],seed[3620],seed[3314],seed[234],seed[3010],seed[486],seed[3554],seed[3278],seed[3711],seed[1818],seed[970],seed[2348],seed[1428],seed[3808],seed[969],seed[881],seed[4094],seed[3841],seed[1662],seed[897],seed[2238],seed[1564],seed[817],seed[4057],seed[2450],seed[1776],seed[3618],seed[3631],seed[2088],seed[3510],seed[1026],seed[1575],seed[4065],seed[72],seed[2696],seed[3801],seed[1568],seed[3566],seed[144],seed[3345],seed[2868],seed[1590],seed[2187],seed[4072],seed[478],seed[3608],seed[1626],seed[590],seed[41],seed[1449],seed[2359],seed[436],seed[442],seed[4089],seed[1630],seed[3192],seed[227],seed[2968],seed[2367],seed[3953],seed[1951],seed[1790],seed[3817],seed[1470],seed[4026],seed[3000],seed[56],seed[2152],seed[1139],seed[2451],seed[3334],seed[2931],seed[3367],seed[190],seed[847],seed[1464],seed[596],seed[862],seed[295],seed[3183],seed[17],seed[832],seed[3464],seed[1527],seed[1393],seed[872],seed[3703],seed[2077],seed[3827],seed[1577],seed[3408],seed[2250],seed[3576],seed[3305],seed[948],seed[773],seed[886],seed[1265],seed[1997],seed[2148],seed[1685],seed[4067],seed[3184],seed[1268],seed[1926],seed[2761],seed[1563],seed[3662],seed[2396],seed[3344],seed[1252],seed[2880],seed[437],seed[1466],seed[627],seed[762],seed[51],seed[842],seed[3293],seed[3068],seed[175],seed[839],seed[1763],seed[1051],seed[3894],seed[1460],seed[149],seed[2157],seed[469],seed[2550],seed[3440],seed[1949],seed[3420],seed[2384],seed[4037],seed[3873],seed[215],seed[1876],seed[2832],seed[357],seed[2374],seed[3571],seed[1090],seed[314],seed[2729],seed[2074],seed[4029],seed[3132],seed[3974],seed[1526],seed[912],seed[529],seed[2944],seed[1326],seed[1089],seed[3394],seed[1827],seed[3306],seed[3995],seed[413],seed[3616],seed[2305],seed[3836],seed[9],seed[4041],seed[1992],seed[1184],seed[3655],seed[2665],seed[1336],seed[2064],seed[3115],seed[81],seed[1586],seed[1272],seed[2200],seed[3418],seed[889],seed[3173],seed[1000],seed[3475],seed[1066],seed[2640],seed[503],seed[2825],seed[2192],seed[1073],seed[3856],seed[2139],seed[1885],seed[2040],seed[254],seed[2821],seed[2167],seed[547],seed[1032],seed[3575],seed[591],seed[2136],seed[1226],seed[3962],seed[1908],seed[471],seed[4068],seed[3357],seed[2205],seed[282],seed[3368],seed[3432],seed[3469],seed[272],seed[2226],seed[180],seed[3990],seed[1160],seed[1037],seed[2062],seed[1679],seed[487],seed[3092],seed[2199],seed[3083],seed[1473],seed[1742],seed[2476],seed[820],seed[1122],seed[3762],seed[217],seed[375],seed[2796],seed[4033],seed[2198],seed[1582],seed[1212],seed[3800],seed[2168],seed[3196],seed[162],seed[2056],seed[1245],seed[2310],seed[4],seed[2259],seed[3866],seed[2309],seed[1389],seed[3329],seed[2302],seed[2470],seed[3997],seed[2497],seed[2789],seed[2731],seed[2611],seed[1003],seed[4022],seed[3426],seed[160],seed[2783],seed[23],seed[2733],seed[1913],seed[3538],seed[2990],seed[3117],seed[3107],seed[537],seed[2381],seed[3710],seed[2453],seed[1502],seed[1723],seed[1384],seed[1772],seed[1902],seed[3333],seed[985],seed[3110],seed[3604],seed[1673],seed[3597],seed[2656],seed[1743],seed[20],seed[1353],seed[1485],seed[3216],seed[1785],seed[3316],seed[1366],seed[693],seed[3546],seed[3875],seed[1102],seed[2882],seed[4011],seed[3019],seed[3986],seed[3633],seed[1260],seed[1831],seed[706],seed[3103],seed[2254],seed[3398],seed[3025],seed[526],seed[3141],seed[3024],seed[3977],seed[2566],seed[3307],seed[1220],seed[826],seed[323],seed[1583],seed[3727],seed[2182],seed[810],seed[1650],seed[224],seed[1321],seed[2142],seed[283],seed[2054],seed[3294],seed[2741],seed[2620],seed[1092],seed[2027],seed[2716],seed[1369],seed[483],seed[715],seed[7],seed[2915],seed[3143],seed[2007],seed[3482],seed[1455],seed[2515],seed[2475],seed[126],seed[990],seed[91],seed[103],seed[992],seed[2176],seed[1532],seed[2045],seed[2456],seed[586],seed[1618],seed[3925],seed[932],seed[3761],seed[3313],seed[1376],seed[1692],seed[3354],seed[2404],seed[1596],seed[755],seed[3382],seed[709],seed[687],seed[2537],seed[3506],seed[2252],seed[2844],seed[1570],seed[580],seed[2746],seed[2117],seed[2145],seed[2684],seed[50],seed[888],seed[100],seed[3422],seed[3343],seed[887],seed[1955],seed[1782],seed[2954],seed[3241],seed[2059],seed[2084],seed[2166],seed[3330],seed[787],seed[3882],seed[3507],seed[1462],seed[1695],seed[523],seed[3553],seed[1192],seed[2999],seed[3412],seed[1415],seed[3219],seed[1423],seed[4056],seed[1099],seed[3876],seed[1283],seed[1198],seed[324],seed[2754],seed[3672],seed[3741],seed[1639],seed[677],seed[1256],seed[3158],seed[2855],seed[3659],seed[770],seed[4063],seed[3171],seed[962],seed[232],seed[2228],seed[1371],seed[55],seed[1029],seed[1234],seed[3541],seed[1698],seed[3119],seed[1886],seed[3347],seed[1629],seed[1825],seed[4082],seed[1615],seed[2337],seed[281],seed[507],seed[3858],seed[570],seed[128],seed[271],seed[1953],seed[3611],seed[430],seed[3522],seed[2560],seed[2745],seed[2097],seed[3750],seed[519],seed[3653],seed[1258],seed[1278],seed[3534],seed[1472],seed[1352],seed[1703],seed[2720],seed[1830],seed[2246],seed[2435],seed[3956],seed[3932],seed[1075],seed[510],seed[216],seed[2350],seed[2235],seed[545],seed[4040],seed[2762],seed[255],seed[3414],seed[1554],seed[2974],seed[276],seed[1900],seed[490],seed[392]}; 
//        seed4 <= {seed[3009],seed[3046],seed[268],seed[200],seed[1455],seed[1031],seed[3307],seed[3096],seed[3119],seed[493],seed[2671],seed[1150],seed[3621],seed[412],seed[3785],seed[2453],seed[2034],seed[3350],seed[3498],seed[3598],seed[2570],seed[3979],seed[1970],seed[902],seed[847],seed[791],seed[1309],seed[404],seed[130],seed[3735],seed[39],seed[1737],seed[3400],seed[3817],seed[3111],seed[2839],seed[3921],seed[3813],seed[3623],seed[1674],seed[3746],seed[4073],seed[483],seed[3831],seed[1110],seed[1806],seed[1384],seed[429],seed[1207],seed[1091],seed[960],seed[749],seed[2389],seed[1360],seed[3195],seed[3468],seed[3728],seed[3044],seed[713],seed[1498],seed[1263],seed[155],seed[3033],seed[3857],seed[3691],seed[1247],seed[1220],seed[2747],seed[3557],seed[1715],seed[562],seed[7],seed[3408],seed[1506],seed[3646],seed[2065],seed[2864],seed[2422],seed[1611],seed[3045],seed[4093],seed[1854],seed[1914],seed[2167],seed[2125],seed[1616],seed[2481],seed[2889],seed[569],seed[4080],seed[2812],seed[987],seed[549],seed[2134],seed[1516],seed[1284],seed[2782],seed[3030],seed[2693],seed[278],seed[1158],seed[3308],seed[3690],seed[3438],seed[3624],seed[2666],seed[2713],seed[1833],seed[1820],seed[2676],seed[12],seed[1633],seed[2658],seed[335],seed[542],seed[2925],seed[1470],seed[3609],seed[574],seed[3645],seed[3605],seed[2896],seed[3680],seed[2630],seed[2610],seed[897],seed[3227],seed[3364],seed[2221],seed[2386],seed[3975],seed[903],seed[2979],seed[3015],seed[3633],seed[3058],seed[2201],seed[399],seed[1156],seed[2659],seed[1035],seed[3446],seed[1074],seed[820],seed[193],seed[3882],seed[3516],seed[3991],seed[1818],seed[2541],seed[2060],seed[666],seed[2727],seed[71],seed[660],seed[3504],seed[3913],seed[99],seed[3283],seed[2072],seed[3812],seed[3767],seed[3532],seed[3346],seed[1234],seed[1959],seed[450],seed[3077],seed[14],seed[1505],seed[3614],seed[1204],seed[817],seed[1072],seed[1011],seed[1965],seed[596],seed[3951],seed[1051],seed[2147],seed[174],seed[2656],seed[804],seed[2959],seed[3215],seed[98],seed[1194],seed[3117],seed[1332],seed[2490],seed[3715],seed[2780],seed[2950],seed[2878],seed[3640],seed[1856],seed[708],seed[3788],seed[3322],seed[2370],seed[1657],seed[1655],seed[838],seed[2249],seed[423],seed[1721],seed[2188],seed[2772],seed[2967],seed[1105],seed[869],seed[3319],seed[2771],seed[4016],seed[2619],seed[711],seed[1858],seed[3896],seed[3368],seed[1756],seed[242],seed[3945],seed[2206],seed[2230],seed[572],seed[3681],seed[2280],seed[181],seed[2284],seed[1160],seed[116],seed[2058],seed[3189],seed[3796],seed[2894],seed[637],seed[754],seed[1282],seed[742],seed[1040],seed[766],seed[1980],seed[2668],seed[2421],seed[3310],seed[2269],seed[59],seed[182],seed[2555],seed[165],seed[682],seed[1705],seed[2022],seed[1998],seed[491],seed[400],seed[720],seed[3964],seed[2568],seed[3130],seed[2567],seed[2688],seed[2363],seed[1610],seed[1813],seed[1411],seed[2311],seed[2182],seed[3049],seed[1169],seed[3328],seed[3843],seed[3141],seed[1971],seed[1672],seed[306],seed[2024],seed[2351],seed[1266],seed[3860],seed[1739],seed[2665],seed[3198],seed[1500],seed[3657],seed[2867],seed[3747],seed[2973],seed[1094],seed[3769],seed[566],seed[1413],seed[2775],seed[2640],seed[3494],seed[3205],seed[1932],seed[3097],seed[593],seed[3886],seed[3524],seed[2598],seed[1210],seed[1696],seed[2604],seed[3210],seed[3039],seed[492],seed[2863],seed[60],seed[1188],seed[1767],seed[1319],seed[3406],seed[3658],seed[4090],seed[2834],seed[2457],seed[1477],seed[2859],seed[272],seed[1046],seed[3148],seed[2492],seed[4060],seed[2231],seed[934],seed[203],seed[1133],seed[2124],seed[967],seed[4046],seed[386],seed[294],seed[2911],seed[845],seed[169],seed[2448],seed[1253],seed[2919],seed[3707],seed[3465],seed[223],seed[1771],seed[1568],seed[3556],seed[2339],seed[1810],seed[1629],seed[2736],seed[420],seed[3334],seed[1566],seed[2843],seed[1837],seed[2399],seed[3485],seed[19],seed[786],seed[3798],seed[725],seed[1957],seed[3125],seed[102],seed[2813],seed[931],seed[3804],seed[1244],seed[1028],seed[3694],seed[1059],seed[3577],seed[1060],seed[2025],seed[119],seed[1324],seed[1826],seed[1708],seed[2765],seed[2857],seed[3288],seed[570],seed[737],seed[1951],seed[2452],seed[3380],seed[1750],seed[3123],seed[115],seed[787],seed[662],seed[2160],seed[878],seed[834],seed[1054],seed[2810],seed[531],seed[1396],seed[263],seed[3133],seed[82],seed[1488],seed[3825],seed[2478],seed[113],seed[597],seed[507],seed[2085],seed[1277],seed[3171],seed[2877],seed[108],seed[2573],seed[776],seed[1988],seed[703],seed[3875],seed[994],seed[2648],seed[2028],seed[2184],seed[3375],seed[527],seed[3251],seed[3729],seed[1982],seed[3292],seed[2396],seed[151],seed[3844],seed[3655],seed[137],seed[3669],seed[1180],seed[627],seed[2788],seed[1582],seed[2687],seed[138],seed[2113],seed[1978],seed[2050],seed[2094],seed[187],seed[1387],seed[831],seed[40],seed[316],seed[1489],seed[3683],seed[3572],seed[112],seed[2618],seed[854],seed[4044],seed[460],seed[1814],seed[362],seed[500],seed[3930],seed[2700],seed[2714],seed[3803],seed[1595],seed[1435],seed[215],seed[2794],seed[1975],seed[674],seed[2491],seed[1699],seed[3137],seed[1613],seed[3032],seed[3037],seed[2070],seed[3706],seed[3667],seed[3642],seed[1353],seed[135],seed[2271],seed[332],seed[2985],seed[1355],seed[1403],seed[1995],seed[396],seed[3026],seed[2746],seed[219],seed[2236],seed[2251],seed[3947],seed[794],seed[1122],seed[31],seed[3588],seed[1786],seed[3933],seed[3379],seed[3267],seed[675],seed[41],seed[3443],seed[1599],seed[545],seed[2850],seed[3279],seed[1717],seed[3779],seed[52],seed[2807],seed[1539],seed[3997],seed[3617],seed[1231],seed[2735],seed[914],seed[1996],seed[3344],seed[3],seed[1223],seed[986],seed[702],seed[2402],seed[663],seed[563],seed[205],seed[1893],seed[2703],seed[2970],seed[671],seed[2243],seed[454],seed[1077],seed[2498],seed[2130],seed[1392],seed[1926],seed[74],seed[1409],seed[1546],seed[3156],seed[3473],seed[1412],seed[3873],seed[1337],seed[3404],seed[3878],seed[1747],seed[1943],seed[3418],seed[2063],seed[315],seed[1710],seed[23],seed[1183],seed[2319],seed[3464],seed[2942],seed[760],seed[4010],seed[2729],seed[2082],seed[1394],seed[941],seed[2428],seed[1153],seed[2384],seed[1646],seed[2446],seed[378],seed[3794],seed[1000],seed[1440],seed[3135],seed[3491],seed[3518],seed[3188],seed[3241],seed[1395],seed[1671],seed[3839],seed[2616],seed[3471],seed[2226],seed[2318],seed[3434],seed[3374],seed[2196],seed[325],seed[3560],seed[1637],seed[937],seed[1200],seed[1476],seed[946],seed[285],seed[2220],seed[2677],seed[624],seed[3367],seed[431],seed[3534],seed[3291],seed[3385],seed[3566],seed[3676],seed[1424],seed[1844],seed[3682],seed[3100],seed[2008],seed[3178],seed[598],seed[107],seed[1534],seed[2509],seed[1731],seed[3483],seed[3738],seed[1380],seed[2081],seed[1149],seed[1103],seed[199],seed[2029],seed[2769],seed[1299],seed[2732],seed[3259],seed[1132],seed[406],seed[3474],seed[1625],seed[1684],seed[3318],seed[976],seed[3731],seed[3153],seed[1903],seed[626],seed[2617],seed[188],seed[680],seed[2635],seed[331],seed[640],seed[829],seed[3463],seed[526],seed[401],seed[2720],seed[3104],seed[2503],seed[1556],seed[1925],seed[3508],seed[1704],seed[437],seed[3819],seed[2836],seed[347],seed[1827],seed[373],seed[345],seed[3601],seed[1983],seed[3360],seed[3711],seed[4089],seed[1084],seed[1316],seed[288],seed[3127],seed[938],seed[573],seed[2062],seed[28],seed[3495],seed[3923],seed[1920],seed[1614],seed[581],seed[2380],seed[1467],seed[745],seed[1656],seed[3401],seed[1673],seed[571],seed[2208],seed[3759],seed[2451],seed[3266],seed[1290],seed[1789],seed[1669],seed[217],seed[1512],seed[2036],seed[2071],seed[1269],seed[1843],seed[51],seed[2104],seed[2033],seed[1991],seed[2506],seed[3685],seed[1466],seed[1388],seed[4088],seed[1815],seed[1691],seed[2578],seed[706],seed[3582],seed[2204],seed[3229],seed[1085],seed[432],seed[2832],seed[3220],seed[3000],seed[1437],seed[158],seed[2296],seed[2507],seed[621],seed[3751],seed[171],seed[2173],seed[2300],seed[3031],seed[2107],seed[2288],seed[1964],seed[2642],seed[1563],seed[1897],seed[1499],seed[783],seed[3602],seed[3632],seed[1314],seed[3353],seed[18],seed[3616],seed[2809],seed[314],seed[3919],seed[1758],seed[3703],seed[3708],seed[2193],seed[1538],seed[2789],seed[1801],seed[4082],seed[2073],seed[2279],seed[1921],seed[81],seed[2026],seed[1723],seed[1013],seed[1587],seed[3166],seed[2934],seed[865],seed[1361],seed[2995],seed[653],seed[2006],seed[2390],seed[1834],seed[3073],seed[899],seed[2234],seed[2624],seed[966],seed[407],seed[2157],seed[66],seed[2023],seed[812],seed[3580],seed[300],seed[380],seed[1985],seed[1639],seed[3720],seed[3845],seed[1586],seed[4064],seed[2368],seed[1227],seed[3496],seed[4071],seed[3705],seed[2653],seed[3349],seed[2487],seed[3074],seed[3576],seed[3355],seed[456],seed[2767],seed[3841],seed[2808],seed[411],seed[1630],seed[616],seed[1064],seed[13],seed[2414],seed[2566],seed[1167],seed[3814],seed[1778],seed[2672],seed[1911],seed[633],seed[9],seed[1176],seed[1181],seed[1930],seed[991],seed[2704],seed[832],seed[3523],seed[2643],seed[3078],seed[1864],seed[1529],seed[3853],seed[1113],seed[2981],seed[2999],seed[2890],seed[789],seed[2185],seed[179],seed[1260],seed[3174],seed[942],seed[1255],seed[2098],seed[2538],seed[1447],seed[308],seed[1627],seed[1137],seed[270],seed[1553],seed[3143],seed[185],seed[3414],seed[2644],seed[3154],seed[2429],seed[2454],seed[814],seed[3028],seed[3884],seed[1984],seed[2365],seed[1608],seed[1565],seed[1313],seed[910],seed[874],seed[2350],seed[3020],seed[591],seed[1386],seed[3990],seed[416],seed[1206],seed[2357],seed[1677],seed[1949],seed[3625],seed[291],seed[2702],seed[2623],seed[1326],seed[45],seed[344],seed[2483],seed[1584],seed[2929],seed[3219],seed[361],seed[3088],seed[2077],seed[235],seed[430],seed[1675],seed[2021],seed[1762],seed[1787],seed[3543],seed[1693],seed[2560],seed[3584],seed[3282],seed[844],seed[143],seed[3050],seed[307],seed[3341],seed[1146],seed[42],seed[3943],seed[1760],seed[2632],seed[3208],seed[3330],seed[722],seed[3949],seed[2508],seed[402],seed[1759],seed[1436],seed[2348],seed[4053],seed[2444],seed[922],seed[908],seed[3458],seed[1378],seed[3663],seed[1623],seed[871],seed[3196],seed[1768],seed[3252],seed[305],seed[3451],seed[3752],seed[1752],seed[2575],seed[2800],seed[1010],seed[3072],seed[2387],seed[2546],seed[1919],seed[2158],seed[718],seed[679],seed[3757],seed[2440],seed[4050],seed[227],seed[3835],seed[781],seed[1119],seed[2456],seed[2980],seed[3678],seed[3739],seed[2937],seed[2759],seed[1907],seed[3548],seed[474],seed[3336],seed[1992],seed[583],seed[1179],seed[3679],seed[417],seed[1860],seed[4079],seed[2493],seed[1873],seed[2106],seed[2138],seed[3014],seed[2516],seed[2057],seed[3022],seed[1067],seed[1532],seed[1274],seed[588],seed[3129],seed[2791],seed[3865],seed[122],seed[1092],seed[1017],seed[2891],seed[3164],seed[958],seed[2885],seed[2069],seed[1257],seed[1915],seed[1159],seed[4014],seed[1305],seed[3562],seed[1716],seed[2627],seed[2056],seed[2340],seed[2172],seed[148],seed[3057],seed[3297],seed[2922],seed[2292],seed[3957],seed[97],seed[128],seed[2753],seed[3052],seed[3412],seed[2673],seed[3920],seed[575],seed[201],seed[1665],seed[520],seed[3699],seed[1405],seed[2913],seed[2792],seed[77],seed[3388],seed[395],seed[2406],seed[144],seed[4028],seed[2531],seed[3828],seed[2449],seed[3898],seed[2411],seed[4055],seed[3615],seed[2636],seed[1558],seed[560],seed[2347],seed[2683],seed[1340],seed[133],seed[2797],seed[732],seed[2997],seed[2593],seed[2317],seed[819],seed[2301],seed[296],seed[3488],seed[1829],seed[3982],seed[2730],seed[3124],seed[534],seed[2032],seed[763],seed[816],seed[1668],seed[1927],seed[2222],seed[1901],seed[3537],seed[3575],seed[1761],seed[289],seed[3186],seed[2198],seed[222],seed[1371],seed[2825],seed[601],seed[777],seed[2191],seed[3940],seed[2875],seed[2265],seed[1987],seed[3815],seed[3163],seed[391],seed[3559],seed[2978],seed[4],seed[2447],seed[72],seed[2123],seed[3637],seed[95],seed[1681],seed[1811],seed[3758],seed[2048],seed[240],seed[3594],seed[2295],seed[2831],seed[2581],seed[3043],seed[2410],seed[3824],seed[2007],seed[1006],seed[1724],seed[2953],seed[2404],seed[3054],seed[1809],seed[2849],seed[343],seed[1358],seed[1288],seed[3326],seed[4002],seed[2290],seed[1391],seed[1254],seed[940],seed[25],seed[2725],seed[644],seed[2115],seed[3021],seed[4067],seed[1297],seed[372],seed[2341],seed[1635],seed[3644],seed[3478],seed[1294],seed[3607],seed[4052],seed[2315],seed[1147],seed[350],seed[4026],seed[3149],seed[2038],seed[2031],seed[780],seed[697],seed[2822],seed[1869],seed[1221],seed[3320],seed[3958],seed[1766],seed[1184],seed[1136],seed[1644],seed[3626],seed[1486],seed[1754],seed[2096],seed[1302],seed[1480],seed[4017],seed[4035],seed[3927],seed[1116],seed[916],seed[1770],seed[2707],seed[1536],seed[1036],seed[3253],seed[1963],seed[3880],seed[2272],seed[3999],seed[1757],seed[2872],seed[694],seed[4062],seed[2554],seed[1725],seed[3959],seed[2010],seed[1073],seed[988],seed[252],seed[2586],seed[3695],seed[3363],seed[2824],seed[1709],seed[1414],seed[2544],seed[3545],seed[1654],seed[1946],seed[3142],seed[1020],seed[1393],seed[1454],seed[2542],seed[1289],seed[2256],seed[959],seed[1268],seed[304],seed[759],seed[79],seed[3549],seed[2382],seed[2883],seed[4038],seed[3387],seed[2171],seed[3005],seed[3883],seed[2267],seed[3087],seed[2726],seed[1124],seed[3976],seed[1853],seed[709],seed[1792],seed[1069],seed[211],seed[3442],seed[3937],seed[2018],seed[394],seed[3131],seed[1492],seed[896],seed[849],seed[214],seed[2868],seed[1323],seed[2461],seed[951],seed[2691],seed[3296],seed[3567],seed[3204],seed[815],seed[1056],seed[3306],seed[1632],seed[62],seed[1478],seed[2227],seed[3822],seed[3132],seed[3324],seed[172],seed[3102],seed[3082],seed[1940],seed[756],seed[194],seed[2881],seed[2907],seed[850],seed[2355],seed[1518],seed[249],seed[2670],seed[3247],seed[837],seed[2304],seed[843],seed[1218],seed[1249],seed[2572],seed[359],seed[3106],seed[3277],seed[2738],seed[298],seed[618],seed[2177],seed[2611],seed[3152],seed[2327],seed[856],seed[3255],seed[1857],seed[3583],seed[2470],seed[700],seed[2874],seed[579],seed[1631],seed[1032],seed[1166],seed[3926],seed[3370],seed[3709],seed[2294],seed[397],seed[836],seed[3238],seed[351],seed[3954],seed[2988],seed[1193],seed[1842],seed[1406],seed[3784],seed[3972],seed[2019],seed[2882],seed[1390],seed[1485],seed[1344],seed[2450],seed[2179],seed[2706],seed[1592],seed[2579],seed[2401],seed[2674],seed[2424],seed[311],seed[891],seed[1976],seed[2375],seed[2865],seed[2485],seed[1428],seed[3659],seed[1471],seed[1561],seed[2212],seed[3864],seed[355],seed[3352],seed[2900],seed[3486],seed[446],seed[1776],seed[1177],seed[568],seed[2861],seed[488],seed[2061],seed[2281],seed[465],seed[2165],seed[654],seed[2606],seed[2285],seed[1140],seed[2298],seed[1900],seed[3335],seed[3967],seed[911],seed[731],seed[2910],seed[164],seed[348],seed[2047],seed[1451],seed[1549],seed[1560],seed[912],seed[150],seed[3953],seed[312],seed[225],seed[243],seed[3487],seed[999],seed[953],seed[1504],seed[747],seed[730],seed[497],seed[1415],seed[3236],seed[3298],seed[1507],seed[2142],seed[3956],seed[2701],seed[75],seed[1062],seed[485],seed[1401],seed[1846],seed[2187],seed[2960],seed[3774],seed[3396],seed[673],seed[717],seed[1431],seed[1003],seed[3382],seed[1913],seed[3521],seed[580],seed[1527],seed[2975],seed[1267],seed[2535],seed[3966],seed[2828],seed[1198],seed[3517],seed[3889],seed[3454],seed[2425],seed[522],seed[161],seed[933],seed[3772],seed[1604],seed[1692],seed[1154],seed[876],seed[3730],seed[3475],seed[2639],seed[641],seed[1531],seed[2823],seed[811],seed[3365],seed[2846],seed[2525],seed[512],seed[3847],seed[3497],seed[3526],seed[1502],seed[2645],seed[585],seed[2592],seed[398],seed[1535],seed[525],seed[3193],seed[603],seed[1670],seed[2122],seed[3392],seed[3946],seed[24],seed[1107],seed[3998],seed[2916],seed[1058],seed[35],seed[748],seed[1803],seed[1589],seed[2600],seed[2977],seed[2009],seed[1548],seed[4015],seed[36],seed[1667],seed[3762],seed[2228],seed[436],seed[2091],seed[689],seed[2126],seed[3460],seed[2499],seed[3608],seed[2376],seed[1005],seed[4083],seed[3978],seed[4030],seed[3915],seed[3677],seed[2553],seed[3323],seed[2286],seed[89],seed[605],seed[1063],seed[1261],seed[2150],seed[1783],seed[1134],seed[2949],seed[602],seed[521],seed[746],seed[3697],seed[1640],seed[3151],seed[2426],seed[3359],seed[1443],seed[247],seed[2246],seed[2373],seed[620],seed[632],seed[455],seed[1609],seed[1322],seed[3611],seed[1519],seed[392],seed[1039],seed[3931],seed[121],seed[617],seed[2833],seed[1753],seed[145],seed[1205],seed[197],seed[2011],seed[1278],seed[1408],seed[178],seed[977],seed[1938],seed[2076],seed[2276],seed[3118],seed[3212],seed[2930],seed[3634],seed[2921],seed[638],seed[1571],seed[297],seed[2099],seed[2948],seed[3013],seed[3453],seed[949],seed[443],seed[2169],seed[303],seed[1969],seed[2958],seed[3895],seed[2408],seed[1429],seed[2001],seed[232],seed[1937],seed[2998],seed[2563],seed[807],seed[1475],seed[1482],seed[3639],seed[1400],seed[2596],seed[2705],seed[890],seed[375],seed[3808],seed[2915],seed[1374],seed[1840],seed[1318],seed[3996],seed[3126],seed[882],seed[950],seed[2074],seed[1093],seed[1583],seed[3300],seed[4074],seed[3613],seed[924],seed[1962],seed[2328],seed[965],seed[3520],seed[3619],seed[3529],seed[2143],seed[3175],seed[1680],seed[228],seed[466],seed[508],seed[2080],seed[2313],seed[2200],seed[650],seed[1125],seed[2356],seed[3936],seed[4004],seed[1083],seed[858],seed[1349],seed[3373],seed[1698],seed[209],seed[3698],seed[3971],seed[1389],seed[2003],seed[3903],seed[1043],seed[3109],seed[3989],seed[2893],seed[2040],seed[2244],seed[505],seed[2178],seed[576],seed[353],seed[3285],seed[2764],seed[91],seed[1356],seed[1808],seed[3112],seed[2161],seed[3480],seed[728],seed[607],seed[4066],seed[1430],seed[3832],seed[3554],seed[1816],seed[2545],seed[652],seed[1828],seed[271],seed[2240],seed[3047],seed[274],seed[3017],seed[2936],seed[1121],seed[877],seed[2684],seed[346],seed[2128],seed[2964],seed[1434],seed[1694],seed[87],seed[424],seed[1591],seed[3356],seed[114],seed[822],seed[1262],seed[2982],seed[1600],seed[2164],seed[3809],seed[4006],seed[1233],seed[3856],seed[913],seed[3775],seed[2361],seed[2739],seed[1372],seed[467],seed[770],seed[1450],seed[2109],seed[3603],seed[661],seed[2966],seed[3377],seed[2250],seed[4047],seed[655],seed[608],seed[1222],seed[969],seed[2842],seed[3648],seed[494],seed[239],seed[909],seed[2030],seed[687],seed[3091],seed[1848],seed[3618],seed[2901],seed[32],seed[715],seed[496],seed[166],seed[926],seed[1228],seed[1805],seed[4091],seed[2420],seed[3984],seed[1933],seed[901],seed[139],seed[830],seed[2749],seed[2170],seed[3098],seed[3718],seed[2695],seed[3362],seed[2622],seed[2441],seed[769],seed[469],seed[2145],seed[2235],seed[801],seed[1474],seed[1928],seed[2879],seed[1765],seed[3421],seed[1178],seed[1835],seed[1420],seed[3834],seed[2612],seed[1590],seed[3675],seed[2757],seed[1606],seed[3952],seed[3278],seed[755],seed[3941],seed[84],seed[1774],seed[963],seed[2273],seed[2131],seed[900],seed[1296],seed[2078],seed[3852],seed[905],seed[1238],seed[1989],seed[2652],seed[1624],seed[1009],seed[2105],seed[490],seed[3234],seed[1023],seed[2924],seed[1544],seed[1034],seed[4007],seed[936],seed[3547],seed[561],seed[3327],seed[3668],seed[1375],seed[4018],seed[69],seed[3888],seed[2268],seed[1952],seed[3505],seed[2391],seed[883],seed[1312],seed[3386],seed[3674],seed[2364],seed[613],seed[471],seed[1866],seed[2946],seed[1095],seed[2751],seed[3622],seed[1821],seed[555],seed[2895],seed[3851],seed[1917],seed[978],seed[1243],seed[805],seed[1330],seed[2067],seed[1979],seed[3961],seed[1345],seed[2603],seed[3411],seed[2637],seed[1799],seed[3413],seed[4000],seed[3258],seed[886],seed[2093],seed[157],seed[1219],seed[948],seed[1252],seed[3546],seed[3665],seed[3743],seed[3929],seed[3912],seed[3908],seed[584],seed[586],seed[125],seed[1785],seed[3140],seed[1459],seed[3760],seed[1742],seed[1626],seed[3745],seed[1923],seed[3089],seed[442],seed[2349],seed[67],seed[2087],seed[3254],seed[2302],seed[1797],seed[2345],seed[3136],seed[1075],seed[1327],seed[1540],seed[635],seed[2761],seed[3818],seed[1550],seed[3450],seed[881],seed[3407],seed[253],seed[1720],seed[2504],seed[3110],seed[301],seed[1385],seed[363],seed[1891],seed[2909],seed[317],seed[547],seed[511],seed[639],seed[2935],seed[3604],seed[1916],seed[2316],seed[1029],seed[3426],seed[772],seed[1446],seed[2260],seed[2321],seed[594],seed[326],seed[3983],seed[3565],seed[3733],seed[729],seed[3850],seed[2785],seed[3969],seed[3416],seed[664],seed[3347],seed[1612],seed[688],seed[2466],seed[3391],seed[3977],seed[3939],seed[3811],seed[1007],seed[3686],seed[379],seed[2016],seed[3980],seed[2951],seed[3402],seed[928],seed[3489],seed[322],seed[2431],seed[767],seed[2395],seed[230],seed[1303],seed[3748],seed[3906],seed[921],seed[221],seed[3661],seed[510],seed[1666],seed[1473],seed[3008],seed[1650],seed[3061],seed[147],seed[3466],seed[458],seed[3372],seed[686],seed[1906],seed[3872],seed[1264],seed[1120],seed[384],seed[3243],seed[2569],seed[1687],seed[866],seed[556],seed[2477],seed[724],seed[980],seed[2550],seed[409],seed[917],seed[3771],seed[1555],seed[2608],seed[1185],seed[589],seed[3034],seed[216],seed[2468],seed[2657],seed[647],seed[2803],seed[1643],seed[2059],seed[2101],seed[1298],seed[2042],seed[3176],seed[3993],seed[1364],seed[971],seed[3717],seed[1607],seed[68],seed[2781],seed[2920],seed[1245],seed[1711],seed[1562],seed[3654],seed[1494],seed[3287],seed[282],seed[1187],seed[1730],seed[309],seed[2561],seed[2799],seed[3786],seed[1577],seed[2841],seed[699],seed[1905],seed[2638],seed[4095],seed[3509],seed[1781],seed[2559],seed[2602],seed[149],seed[117],seed[1004],seed[3740],seed[3535],seed[2941],seed[1367],seed[1572],seed[788],seed[1291],seed[1664],seed[302],seed[930],seed[207],seed[751],seed[1130],seed[719],seed[2479],seed[3606],seed[1888],seed[3250],seed[1745],seed[2181],seed[1129],seed[3085],seed[275],seed[2218],seed[735],seed[1131],seed[2917],seed[3261],seed[4022],seed[390],seed[1918],seed[1163],seed[109],seed[448],seed[3826],seed[2151],seed[2027],seed[90],seed[3536],seed[2938],seed[1143],seed[3122],seed[377],seed[543],seed[495],seed[1079],seed[3628],seed[472],seed[177],seed[1071],seed[3684],seed[3120],seed[1875],seed[1172],seed[3514],seed[3165],seed[2084],seed[875],seed[3948],seed[3286],seed[3573],seed[4057],seed[356],seed[4019],seed[3909],seed[504],seed[3827],seed[1295],seed[57],seed[860],seed[3419],seed[3209],seed[2360],seed[3029],seed[3477],seed[4008],seed[1567],seed[170],seed[3002],seed[2342],seed[2562],seed[58],seed[1662],seed[3482],seed[2811],seed[984],seed[3519],seed[3224],seed[2472],seed[393],seed[428],seed[3035],seed[3256],seed[2183],seed[2203],seed[2053],seed[2320],seed[3274],seed[611],seed[658],seed[2523],seed[710],seed[1645],seed[2412],seed[3312],seed[3228],seed[2745],seed[1369],seed[1794],seed[281],seed[2871],seed[1986],seed[3018],seed[2821],seed[1545],seed[774],seed[4020],seed[3260],seed[636],seed[1037],seed[1763],seed[2192],seed[907],seed[2862],seed[544],seed[761],seed[2718],seed[1239],seed[1022],seed[4045],seed[2679],seed[2983],seed[1523],seed[2002],seed[3108],seed[3447],seed[3113],seed[3636],seed[3599],seed[993],seed[1108],seed[3870],seed[123],seed[2787],seed[3430],seed[167],seed[1735],seed[532],seed[3290],seed[3492],seed[146],seed[683],seed[892],seed[2486],seed[919],seed[685],seed[2912],seed[2888],seed[3742],seed[1270],seed[1772],seed[2464],seed[3284],seed[990],seed[2796],seed[1283],seed[1881],seed[1990],seed[2004],seed[389],seed[1524],seed[105],seed[1216],seed[1647],seed[853],seed[3476],seed[2136],seed[1511],seed[3202],seed[1841],seed[1484],seed[1383],seed[3107],seed[813],seed[1559],seed[3265],seed[435],seed[3099],seed[3422],seed[2918],seed[1338],seed[295],seed[1379],seed[3144],seed[524],seed[3805],seed[2664],seed[1968],seed[3182],seed[2969],seed[1065],seed[2584],seed[2580],seed[3056],seed[1462],seed[894],seed[1936],seed[3836],seed[1569],seed[2309],seed[1086],seed[3019],seed[4025],seed[425],seed[3833],seed[2906],seed[365],seed[2991],seed[3539],seed[1135],seed[2518],seed[1885],seed[1743],seed[1839],seed[2369],seed[864],seed[2520],seed[3242],seed[1448],seed[56],seed[333],seed[4043],seed[76],seed[83],seed[1780],seed[352],seed[3838],seed[2416],seed[369],seed[1317],seed[1142],seed[2766],seed[3462],seed[806],seed[2529],seed[3369],seed[37],seed[3907],seed[2536],seed[3868],seed[590],seed[2710],seed[2495],seed[1495],seed[2140],seed[2721],seed[3249],seed[3592],seed[2892],seed[2549],seed[357],seed[3595],seed[2116],seed[3849],seed[4078],seed[3354],seed[3399],seed[3079],seed[3395],seed[1934],seed[1170],seed[476],seed[3167],seed[2014],seed[2335],seed[3631],seed[600],seed[2540],seed[762],seed[3701],seed[2628],seed[1080],seed[478],seed[3922],seed[995],seed[1491],seed[3281],seed[553],seed[403],seed[127],seed[2275],seed[142],seed[364],seed[557],seed[3656],seed[2931],seed[3301],seed[3424],seed[3345],seed[2257],seed[773],seed[4012],seed[2174],seed[3068],seed[669],seed[1580],seed[3459],seed[163],seed[2409],seed[2278],seed[1777],seed[175],seed[2020],seed[3276],seed[2205],seed[3714],seed[3332],seed[3670],seed[1890],seed[2692],seed[1802],seed[463],seed[1877],seed[1878],seed[1701],seed[1859],seed[3435],seed[800],seed[1751],seed[3507],seed[3778],seed[4054],seed[2770],seed[1678],seed[1953],seed[1088],seed[224],seed[1728],seed[93],seed[3510],seed[970],seed[943],seed[1960],seed[3861],seed[2144],seed[3791],seed[2698],seed[798],seed[1224],seed[1514],seed[2066],seed[1686],seed[552],seed[3724],seed[3134],seed[867],seed[3420],seed[3935],seed[989],seed[3837],seed[64],seed[3007],seed[1],seed[529],seed[3425],seed[1882],seed[1196],seed[1898],seed[1068],seed[33],seed[4001],seed[2744],seed[2972],seed[444],seed[3540],seed[1444],seed[604],seed[1237],seed[1399],seed[2697],seed[2459],seed[1024],seed[3070],seed[1453],seed[3036],seed[3799],seed[173],seed[3763],seed[1557],seed[1419],seed[1570],seed[427],seed[1576],seed[2858],seed[1346],seed[2049],seed[3173],seed[2957],seed[473],seed[3503],seed[1706],seed[1526],seed[2869],seed[1033],seed[3066],seed[1427],seed[2838],seed[2168],seed[3076],seed[3965],seed[1300],seed[141],seed[741],seed[481],seed[2211],seed[2681],seed[3862],seed[1879],seed[3216],seed[2620],seed[1530],seed[2835],seed[514],seed[3893],seed[1733],seed[1061],seed[523],seed[2287],seed[1273],seed[2141],seed[872],seed[1804],seed[707],seed[3741],seed[2576],seed[2075],seed[1001],seed[2255],seed[2994],seed[2176],seed[382],seed[2088],seed[1100],seed[828],seed[233],seed[4092],seed[1329],seed[176],seed[550],seed[1041],seed[810],seed[4068],seed[2898],seed[3423],seed[2526],seed[2962],seed[1162],seed[1966],seed[3973],seed[383],seed[1588],seed[2366],seed[3689],seed[261],seed[785],seed[3859],seed[3147],seed[1552],seed[3571],seed[595],seed[1026],seed[238],seed[3321],seed[3866],seed[3924],seed[2961],seed[2565],seed[3820],seed[1605],seed[2927],seed[2945],seed[3063],seed[3635],seed[721],seed[3773],seed[964],seed[665],seed[236],seed[3754],seed[2139],seed[499],seed[2473],seed[2851],seed[2552],seed[968],seed[2837],seed[1830],seed[2442],seed[1522],seed[132],seed[1214],seed[3191],seed[1967],seed[1164],seed[2774],seed[2352],seed[1973],seed[1173],seed[2153],seed[503],seed[939],seed[3311],seed[2845],seed[2371],seed[3515],seed[3855],seed[2397],seed[1417],seed[3275],seed[3499],seed[4048],seed[578],seed[1543],seed[740],seed[873],seed[1999],seed[2166],seed[2805],seed[1025],seed[323],seed[3337],seed[3702],seed[645],seed[2467],seed[2407],seed[2820],seed[577],seed[1542],seed[3810],seed[2990],seed[461],seed[1321],seed[1398],seed[1904],seed[2312],seed[2334],seed[3552],seed[2114],seed[3449],seed[516],seed[2329],seed[2660],seed[3168],seed[256],seed[1203],seed[2795],seed[506],seed[276],seed[3159],seed[2133],seed[3180],seed[1320],seed[2694],seed[1141],seed[2358],seed[2923],seed[3790],seed[1547],seed[2776],seed[3721],seed[3673],seed[3272],seed[370],seed[3610],seed[1148],seed[2615],seed[2699],seed[2758],seed[3726],seed[3158],seed[753],seed[1910],seed[3383],seed[1867],seed[2500],seed[2484],seed[1902],seed[2353],seed[4084],seed[1157],seed[539],seed[3394],seed[3649],seed[3666],seed[3389],seed[3985],seed[733],seed[1045],seed[21],seed[2582],seed[2223],seed[3522],seed[1714],seed[3366],seed[1225],seed[106],seed[935],seed[1748],seed[1537],seed[2354],seed[1793],seed[1248],seed[3011],seed[381],seed[1950],seed[861],seed[3217],seed[1883],seed[691],seed[839],seed[1190],seed[3848],seed[1689],seed[1191],seed[2388],seed[1690],seed[3693],seed[3479],seed[484],seed[3440],seed[3439],seed[3351],seed[1497],seed[2965],seed[559],seed[1510],seed[2992],seed[2336],seed[3986],seed[1702],seed[1382],seed[1886],seed[1469],seed[3218],seed[1452],seed[2557],seed[1870],seed[833],seed[1594],seed[482],seed[1445],seed[2344],seed[2310],seed[2045],seed[2512],seed[1307],seed[771],seed[3995],seed[1246],seed[2064],seed[3981],seed[796],seed[3713],seed[2571],seed[2621],seed[1769],seed[2590],seed[3876],seed[541],seed[868],seed[1070],seed[2149],seed[2847],seed[643],seed[4034],seed[2855],seed[1663],seed[3761],seed[3264],seed[318],seed[254],seed[213],seed[3358],seed[2476],seed[3725],seed[3787],seed[3511],seed[1211],seed[290],seed[3190],seed[489],seed[3756],seed[1880],seed[3145],seed[1659],seed[3512],seed[2806],seed[623],seed[592],seed[3172],seed[1117],seed[3581],seed[3436],seed[6],seed[1128],seed[2000],seed[3867],seed[2475],seed[2417],seed[3452],seed[2213],seed[2238],seed[1351],seed[3177],seed[915],seed[3333],seed[793],seed[587],seed[1603],seed[328],seed[2986],seed[1433],seed[1139],seed[1528],seed[2362],seed[957],seed[1501],seed[634],seed[3080],seed[1597],seed[2902],seed[1838],seed[2784],seed[20],seed[1865],seed[954],seed[548],seed[3716],seed[2303],seed[2588],seed[2634],seed[3115],seed[4013],seed[299],seed[2914],seed[4027],seed[1242],seed[2625],seed[3968],seed[2186],seed[2741],seed[479],seed[765],seed[1740],seed[1638],seed[2458],seed[1513],seed[1106],seed[648],seed[752],seed[3304],seed[3643],seed[2731],seed[2293],seed[1764],seed[1948],seed[2513],seed[2239],seed[2330],seed[3987],seed[3470],seed[1945],seed[3938],seed[2299],seed[2530],seed[1483],seed[1016],seed[2963],seed[2259],seed[1695],seed[4085],seed[1310],seed[2005],seed[3586],seed[1301],seed[2393],seed[893],seed[3071],seed[3789],seed[1863],seed[3890],seed[678],seed[744],seed[186],seed[319],seed[2323],seed[248],seed[2740],seed[120],seed[2403],seed[1642],seed[1636],seed[2155],seed[53],seed[73],seed[4041],seed[2097],seed[321],seed[540],seed[3003],seed[2651],seed[2844],seed[629],seed[2118],seed[2261],seed[809],seed[681],seed[1050],seed[895],seed[2607],seed[180],seed[2522],seed[29],seed[2750],seed[1335],seed[714],seed[3877],seed[2534],seed[63],seed[985],seed[818],seed[422],seed[3398],seed[2089],seed[2870],seed[2055],seed[1165],seed[3472],seed[3513],seed[1700],seed[1442],seed[3871],seed[3710],seed[1736],seed[842],seed[1896],seed[1352],seed[3530],seed[3232],seed[2111],seed[360],seed[3161],seed[823],seed[3630],seed[3490],seed[2194],seed[27],seed[509],seed[2180],seed[857],seed[367],seed[1574],seed[2214],seed[4058],seed[3842],seed[615],seed[1517],seed[3469],seed[3139],seed[1463],seed[2886],seed[2337],seed[1258],seed[3315],seed[136],seed[153],seed[2626],seed[1030],seed[1272],seed[2480],seed[313],seed[2463],seed[204],seed[565],seed[2829],seed[2742],seed[1076],seed[3591],seed[3361],seed[1874],seed[3160],seed[2283],seed[3647],seed[3455],seed[3213],seed[2306],seed[2678],seed[3092],seed[2777],seed[631],seed[96],seed[3342],seed[2162],seed[1441],seed[1012],seed[86],seed[2722],seed[341],seed[1791],seed[4003],seed[2215],seed[3750],seed[981],seed[162],seed[1087],seed[2209],seed[3900],seed[925],seed[55],seed[3528],seed[764],seed[3138],seed[649],seed[2202],seed[3331],seed[3223],seed[2233],seed[3025],seed[1350],seed[212],seed[2224],seed[2217],seed[3075],seed[2779],seed[2908],seed[258],seed[3257],seed[2394],seed[1311],seed[1726],seed[3294],seed[3340],seed[1872],seed[3114],seed[1641],seed[3121],seed[1306],seed[2716],seed[3846],seed[220],seed[2591],seed[269],seed[1954],seed[2496],seed[1653],seed[1357],seed[1048],seed[152],seed[3157],seed[1851],seed[2443],seed[3578],seed[1620],seed[2433],seed[1541],seed[808],seed[2826],seed[1651],seed[457],seed[3429],seed[2083],seed[2989],seed[2984],seed[1795],seed[234],seed[1402],seed[3650],seed[1199],seed[2754],seed[1850],seed[1334],seed[1718],seed[4024],seed[3185],seed[3879],seed[889],seed[1102],seed[50],seed[1515],seed[1734],seed[502],seed[3916],seed[651],seed[449],seed[3770],seed[974],seed[2262],seed[464],seed[1852],seed[982],seed[293],seed[3776],seed[513],seed[3950],seed[339],seed[26],seed[3764],seed[3244],seed[2786],seed[1573],seed[3736],seed[2932],seed[1676],seed[3963],seed[2482],seed[5],seed[3461],seed[1280],seed[1057],seed[3894],seed[2551],seed[736],seed[245],seed[3197],seed[2712],seed[3887],seed[1941],seed[920],seed[2926],seed[2996],seed[2884],seed[3280],seed[480],seed[528],seed[1712],seed[2737],seed[1683],seed[992],seed[698],seed[1397],seed[3732],seed[705],seed[3427],seed[1741],seed[354],seed[2241],seed[1575],seed[2680],seed[78],seed[2947],seed[3830],seed[2816],seed[2419],seed[1823],seed[3579],seed[2343],seed[3585],seed[2675],seed[3590],seed[515],seed[3187],seed[3060],seed[4009],seed[3942],seed[3840],seed[3806],seed[47],seed[30],seed[668],seed[3538],seed[3816],seed[716],seed[4086],seed[2135],seed[1285],seed[2514],seed[609],seed[2956],seed[3006],seed[1027],seed[184],seed[2519],seed[1363],seed[690],seed[419],seed[410],seed[2631],seed[599],seed[1449],seed[1053],seed[1021],seed[2210],seed[2661],seed[1884],seed[1275],seed[3671],seed[961],seed[100],seed[551],seed[3672],seed[4069],seed[3795],seed[104],seed[2528],seed[2646],seed[3230],seed[1822],seed[2120],seed[447],seed[2663],seed[468],seed[3417],seed[3203],seed[2974],seed[803],seed[438],seed[61],seed[3874],seed[3542],seed[2558],seed[1145],seed[1496],seed[955],seed[3444],seed[3569],seed[537],seed[462],seed[1460],seed[1118],seed[4056],seed[2719],seed[43],seed[2325],seed[2225],seed[619],seed[1215],seed[168],seed[3829],seed[2943],seed[2359],seed[3660],seed[1832],seed[3782],seed[3823],seed[3574],seed[1719],seed[415],seed[2367],seed[445],seed[704],seed[3181],seed[1015],seed[3206],seed[3289],seed[1368],seed[260],seed[3651],seed[3988],seed[34],seed[2346],seed[945],seed[190],seed[3905],seed[672],seed[3371],seed[3551],seed[3105],seed[997],seed[2815],seed[126],seed[3629],seed[998],seed[1425],seed[198],seed[2372],seed[2728],seed[3314],seed[3313],seed[1790],seed[3027],seed[973],seed[3090],seed[567],seed[2599],seed[797],seed[1189],seed[4077],seed[237],seed[726],seed[2052],seed[2733],seed[784],seed[1161],seed[1342],seed[3722],seed[1333],seed[241],seed[642],seed[1339],seed[2331],seed[2587],seed[2054],seed[1341],seed[1479],seed[1564],seed[1824],seed[2955],seed[3558],seed[2801],seed[2044],seed[3653],seed[202],seed[286],seed[3271],seed[3221],seed[3214],seed[1049],seed[790],seed[310],seed[1366],seed[3299],seed[2445],seed[3664],seed[1648],seed[3184],seed[2515],seed[1315],seed[2253],seed[349],seed[196],seed[231],seed[2987],seed[3792],seed[3409],seed[1018],seed[2497],seed[3700],seed[3723],seed[2667],seed[3970],seed[3914],seed[3169],seed[1410],seed[44],seed[2307],seed[927],seed[646],seed[558],seed[70],seed[1956],seed[3194],seed[336],seed[340],seed[368],seed[1707],seed[4065],seed[2189],seed[3777],seed[1055],seed[2086],seed[3245],seed[743],seed[2148],seed[3428],seed[792],seed[4011],seed[284],seed[3051],seed[1722],seed[2041],seed[1287],seed[944],seed[1362],seed[262],seed[2669],seed[1652],seed[3753],seed[1328],seed[2494],seed[622],seed[1168],seed[3086],seed[779],seed[2804],seed[2852],seed[1197],seed[879],seed[2933],seed[2903],seed[110],seed[1847],seed[782],seed[1876],seed[3305],seed[1598],seed[1418],seed[1426],seed[2332],seed[3231],seed[2108],seed[3917],seed[4031],seed[1658],seed[1939],seed[3962],seed[477],seed[11],seed[2853],seed[1127],seed[2471],seed[434],seed[1174],seed[852],seed[1308],seed[388],seed[1798],seed[582],seed[712],seed[49],seed[696],seed[3235],seed[1082],seed[3433],seed[3162],seed[1861],seed[366],seed[3881],seed[2944],seed[2517],seed[501],seed[3620],seed[244],seed[3128],seed[2110],seed[1871],seed[2489],seed[3555],seed[2079],seed[3593],seed[1279],seed[3596],seed[3493],seed[3042],seed[3797],seed[2474],seed[1042],seed[1679],seed[1421],seed[888],seed[2887],seed[2199],seed[3899],seed[4029],seed[3239],seed[1922],seed[3918],seed[2501],seed[1912],seed[475],seed[887],seed[3587],seed[208],seed[1464],seed[2095],seed[2717],seed[1908],seed[2734],seed[2232],seed[2434],seed[2015],seed[2381],seed[1775],seed[433],seed[1729],seed[2308],seed[3734],seed[3925],seed[3317],seed[4021],seed[947],seed[374],seed[1354],seed[3378],seed[2430],seed[2314],seed[606],seed[183],seed[1038],seed[1099],seed[80],seed[1782],seed[3329],seed[996],seed[2830],seed[2521],seed[2400],seed[3293],seed[2601],seed[870],seed[1457],seed[3041],seed[3527],seed[2511],seed[2068],seed[2121],seed[2564],seed[1807],seed[3016],seed[802],seed[3083],seed[1458],seed[279],seed[2899],seed[693],seed[2305],seed[452],seed[848],seed[3376],seed[3597],seed[3544],seed[824],seed[1104],seed[218],seed[1812],seed[1438],seed[2585],seed[16],seed[1487],seed[2876],seed[1195],seed[1800],seed[1212],seed[1202],seed[265],seed[1098],seed[3944],seed[255],seed[684],seed[1493],seed[3055],seed[3397],seed[2297],seed[1788],seed[4051],seed[266],seed[1240],seed[1688],seed[1944],seed[3854],seed[440],seed[2860],seed[342],seed[2438],seed[2469],seed[376],seed[2012],seed[1052],seed[1713],seed[134],seed[1256],seed[906],seed[2439],seed[414],seed[1836],seed[904],seed[3719],seed[3010],seed[2539],seed[1602],seed[2589],seed[3316],seed[1993],seed[2460],seed[160],seed[2405],seed[3807],seed[3343],seed[3065],seed[564],seed[1596],seed[250],seed[103],seed[2242],seed[1423],seed[4023],seed[2190],seed[264],seed[3116],seed[1336],seed[1490],seed[486],seed[2247],seed[453],seed[2156],seed[825],seed[2817],seed[1579],seed[1090],seed[2819],seed[2119],seed[3688],seed[846],seed[3793],seed[3869],seed[3155],seed[4040],seed[3652],seed[3897],seed[283],seed[3910],seed[2873],seed[3783],seed[3765],seed[821],seed[1465],seed[2723],seed[3103],seed[3589],seed[962],seed[2037],seed[2413],seed[1732],seed[2708],seed[1855],seed[3766],seed[2132],seed[3934],seed[15],seed[1373],seed[2435],seed[3390],seed[3568],seed[1276],seed[3338],seed[1585],seed[533],seed[3641],seed[1554],seed[1407],seed[320],seed[470],seed[835],seed[1619],seed[1892],seed[3393],seed[3309],seed[3062],seed[2848],seed[3432],seed[3038],seed[3094],seed[2270],seed[1796],seed[3437],seed[3211],seed[2755],seed[4087],seed[1370],seed[1304],seed[676],seed[1601],seed[3932],seed[851],seed[3457],seed[1503],seed[3384],seed[3325],seed[3863],seed[3467],seed[48],seed[1123],seed[94],seed[1432],seed[267],seed[54],seed[1002],seed[2709],seed[1192],seed[3911],seed[2129],seed[884],seed[1685],seed[2854],seed[795],seed[4049],seed[2940],seed[2],seed[2046],seed[739],seed[2462],seed[929],seed[3248],seed[1909],seed[206],seed[3500],seed[1365],seed[2245],seed[2374],seed[2103],seed[1481],seed[330],seed[2277],seed[2207],seed[1935],seed[1744],seed[3502],seed[4075],seed[2533],seed[3901],seed[3561],seed[3892],seed[2465],seed[2715],seed[2100],seed[1825],seed[695],seed[841],seed[3994],seed[3273],seed[2237],seed[2548],seed[826],seed[426],seed[3506],seed[1520],seed[1209],seed[692],seed[1622],seed[1784],seed[3403],seed[2197],seed[2968],seed[277],seed[1887],seed[2798],seed[727],seed[1089],seed[2952],seed[3445],seed[3712],seed[2195],seed[1618],seed[2527],seed[2605],seed[3012],seed[88],seed[498],seed[3550],seed[2743],seed[614],seed[1862],seed[3687],seed[385],seed[2971],seed[2383],seed[1376],seed[3339],seed[677],seed[2043],seed[2432],seed[898],seed[657],seed[2633],seed[2609],seed[1931],seed[3612],seed[3501],seed[2013],seed[1292],seed[2017],seed[2090],seed[287],seed[3902],seed[3170],seed[1096],seed[2415],seed[1241],seed[3410],seed[1151],seed[1660],seed[3441],seed[610],seed[1593],seed[273],seed[778],seed[1155],seed[4037],seed[2939],seed[3553],seed[538],seed[2333],seed[750],seed[3246],seed[2595],seed[131],seed[2597],seed[101],seed[2254],seed[1271],seed[3456],seed[1232],seed[554],seed[2904],seed[3415],seed[1894],seed[2928],seed[862],seed[1779],seed[2641],seed[2790],seed[3563],seed[4063],seed[2524],seed[775],seed[2724],seed[1581],seed[118],seed[3302],seed[1578],seed[1738],seed[2127],seed[2175],seed[956],seed[612],seed[1044],seed[226],seed[2686],seed[1889],seed[1929],seed[1994],seed[2897],seed[2488],seed[3801],seed[1727],seed[2654],seed[459],seed[2577],seed[2117],seed[1152],seed[1138],seed[191],seed[1617],seed[1439],seed[3802],seed[3600],seed[111],seed[517],seed[10],seed[1381],seed[1325],seed[1182],seed[3192],seed[2092],seed[3885],seed[1008],seed[2137],seed[880],seed[3295],seed[923],seed[2655],seed[701],seed[1509],seed[863],seed[1097],seed[1817],seed[2154],seed[3448],seed[1236],seed[3781],seed[3744],seed[2556],seed[4081],seed[257],seed[2840],seed[2814],seed[3023],seed[3800],seed[1286],seed[1175],seed[4033],seed[546],seed[4039],seed[2248],seed[3960],seed[3233],seed[3533],seed[2802],seed[3150],seed[979],seed[1468],seed[670],seed[734],seed[154],seed[983],seed[1422],seed[3207],seed[1109],seed[1819],seed[1019],seed[1416],seed[1746],seed[3269],seed[2762],seed[1259],seed[2685],seed[1229],seed[1942],seed[441],seed[3225],seed[2993],seed[2377],seed[2690],seed[1014],seed[439],seed[2282],seed[2035],seed[192],seed[1348],seed[3357],seed[535],seed[3268],seed[799],seed[2326],seed[1961],seed[1217],seed[259],seed[2711],seed[3200],seed[3179],seed[2418],seed[2219],seed[4072],seed[3431],seed[2146],seed[2818],seed[4032],seed[3780],seed[292],seed[1697],seed[1078],seed[2510],seed[334],seed[22],seed[1749],seed[738],seed[1661],seed[2954],seed[3692],seed[3904],seed[3263],seed[518],seed[4036],seed[3992],seed[2427],seed[1955],seed[3262],seed[2266],seed[2437],seed[2547],seed[2905],seed[2662],seed[129],seed[3048],seed[3064],seed[413],seed[2423],seed[2689],seed[1213],seed[3040],seed[4042],seed[2112],seed[4005],seed[3704],seed[2696],seed[1525],seed[2682],seed[3084],seed[3858],seed[1972],seed[1171],seed[4076],seed[2378],seed[1101],seed[2385],seed[2760],seed[3737],seed[1343],seed[0],seed[3237],seed[1226],seed[2436],seed[2264],seed[1924],seed[2793],seed[2159],seed[2614],seed[2102],seed[2051],seed[3541],seed[1251],seed[92],seed[17],seed[952],seed[1112],seed[1533],seed[327],seed[3727],seed[758],seed[2039],seed[1773],seed[2229],seed[3525],seed[3146],seed[1958],seed[3001],seed[975],seed[3570],seed[4070],seed[246],seed[1551],seed[859],seed[210],seed[3755],seed[2322],seed[1461],seed[3696],seed[4061],seed[1230],seed[1845],seed[1456],seed[536],seed[371],seed[2392],seed[1377],seed[3481],seed[530],seed[195],seed[280],seed[2763],seed[656],seed[2752],seed[1281],seed[2613],seed[4094],seed[1628],seed[1521],seed[156],seed[338],seed[3270],seed[2543],seed[1081],seed[1755],seed[3201],seed[3183],seed[2263],seed[2866],seed[3821],seed[2291],seed[2649],seed[1115],seed[2398],seed[2574],seed[855],seed[2502],seed[768],seed[1981],seed[124],seed[2252],seed[2532],seed[1066],seed[1404],seed[1201],seed[329],seed[1186],seed[2505],seed[2778],seed[3627],seed[2583],seed[2768],seed[1974],seed[487],seed[630],seed[2748],seed[2594],seed[408],seed[140],seed[1634],seed[3749],seed[1114],seed[1359],seed[324],seed[159],seed[3101],seed[659],seed[2258],seed[1331],seed[2856],seed[3222],seed[1849],seed[3303],seed[1947],seed[1621],seed[2338],seed[85],seed[840],seed[932],seed[1868],seed[2650],seed[358],seed[827],seed[1144],seed[1977],seed[3891],seed[3564],seed[625],seed[4059],seed[2629],seed[1111],seed[2324],seed[1895],seed[2379],seed[3974],seed[1508],seed[229],seed[628],seed[38],seed[3531],seed[2756],seed[1703],seed[387],seed[1126],seed[1899],seed[3081],seed[2289],seed[2216],seed[8],seed[1997],seed[3067],seed[2773],seed[3004],seed[3348],seed[421],seed[1682],seed[3405],seed[3928],seed[405],seed[757],seed[3662],seed[189],seed[723],seed[3059],seed[65],seed[1649],seed[2455],seed[1250],seed[1347],seed[1265],seed[2976],seed[3768],seed[2163],seed[3053],seed[3199],seed[667],seed[3095],seed[418],seed[1293],seed[337],seed[1472],seed[2880],seed[3638],seed[1208],seed[2274],seed[519],seed[3381],seed[3069],seed[3226],seed[3484],seed[2783],seed[885],seed[1235],seed[972],seed[3024],seed[1047],seed[3240],seed[2647],seed[1615],seed[3955],seed[46],seed[2537],seed[251],seed[2152],seed[451],seed[1831],seed[3093],seed[918],seed[2827]}; 
//        seed5 <= {seed[2337],seed[1934],seed[1406],seed[2097],seed[1209],seed[623],seed[2156],seed[2843],seed[3321],seed[2529],seed[1042],seed[617],seed[227],seed[636],seed[2499],seed[2679],seed[396],seed[882],seed[2662],seed[3776],seed[3946],seed[3628],seed[1082],seed[3061],seed[1675],seed[3639],seed[2907],seed[990],seed[2563],seed[3837],seed[1030],seed[3616],seed[3144],seed[1670],seed[2038],seed[2865],seed[2167],seed[3093],seed[3733],seed[3081],seed[1625],seed[3676],seed[3025],seed[3454],seed[484],seed[3100],seed[2113],seed[1129],seed[715],seed[3045],seed[1328],seed[1038],seed[2225],seed[2164],seed[3929],seed[3147],seed[1172],seed[945],seed[3720],seed[1390],seed[278],seed[3356],seed[3878],seed[651],seed[3413],seed[933],seed[1352],seed[3752],seed[3692],seed[2240],seed[2789],seed[112],seed[1431],seed[3654],seed[2596],seed[621],seed[2311],seed[3652],seed[2218],seed[2883],seed[3274],seed[1252],seed[2964],seed[2166],seed[1800],seed[372],seed[2356],seed[521],seed[3175],seed[3912],seed[4022],seed[1037],seed[2944],seed[3255],seed[2953],seed[1467],seed[2176],seed[2556],seed[1768],seed[1512],seed[3031],seed[123],seed[837],seed[3779],seed[1210],seed[902],seed[2895],seed[1391],seed[738],seed[2109],seed[1114],seed[821],seed[1147],seed[2458],seed[972],seed[1740],seed[3816],seed[3780],seed[2009],seed[3207],seed[813],seed[81],seed[644],seed[1191],seed[1382],seed[3458],seed[1417],seed[3542],seed[3861],seed[1557],seed[3462],seed[1614],seed[3990],seed[1872],seed[3782],seed[2005],seed[3334],seed[1330],seed[384],seed[3104],seed[4063],seed[734],seed[3787],seed[512],seed[3243],seed[2608],seed[1908],seed[2383],seed[1485],seed[236],seed[53],seed[1696],seed[576],seed[2373],seed[1663],seed[1763],seed[3727],seed[1664],seed[1769],seed[452],seed[113],seed[2721],seed[3027],seed[13],seed[3544],seed[3532],seed[3993],seed[1795],seed[3171],seed[3739],seed[3295],seed[2191],seed[539],seed[2532],seed[2574],seed[3710],seed[2346],seed[475],seed[2763],seed[489],seed[3869],seed[1111],seed[591],seed[2654],seed[72],seed[733],seed[300],seed[1651],seed[3392],seed[936],seed[2619],seed[987],seed[662],seed[2444],seed[3037],seed[1597],seed[3564],seed[2023],seed[3914],seed[1883],seed[420],seed[3693],seed[1238],seed[947],seed[3264],seed[2727],seed[4046],seed[2677],seed[3999],seed[811],seed[1929],seed[3862],seed[3822],seed[3437],seed[2012],seed[1548],seed[2811],seed[2650],seed[1452],seed[1949],seed[3279],seed[1353],seed[2448],seed[3358],seed[3699],seed[1764],seed[2273],seed[732],seed[2836],seed[2110],seed[30],seed[391],seed[1882],seed[3096],seed[1412],seed[3698],seed[3103],seed[1376],seed[2316],seed[216],seed[96],seed[2745],seed[142],seed[602],seed[2586],seed[2561],seed[1277],seed[307],seed[3870],seed[3026],seed[3823],seed[2548],seed[2293],seed[2613],seed[1263],seed[2967],seed[3339],seed[741],seed[1011],seed[3820],seed[3346],seed[2050],seed[543],seed[2656],seed[1954],seed[1781],seed[3051],seed[41],seed[2],seed[831],seed[11],seed[3700],seed[3677],seed[1013],seed[1043],seed[2090],seed[509],seed[347],seed[2894],seed[2011],seed[2231],seed[2801],seed[3411],seed[1688],seed[1427],seed[867],seed[298],seed[3706],seed[725],seed[329],seed[1257],seed[1531],seed[373],seed[3017],seed[1225],seed[1092],seed[1824],seed[706],seed[542],seed[2436],seed[27],seed[736],seed[879],seed[392],seed[2220],seed[1308],seed[2179],seed[1091],seed[2234],seed[1870],seed[3962],seed[2454],seed[1451],seed[2208],seed[1957],seed[3432],seed[3245],seed[1060],seed[3858],seed[1588],seed[2777],seed[1628],seed[1029],seed[3211],seed[1283],seed[150],seed[1141],seed[4059],seed[3079],seed[116],seed[845],seed[1259],seed[3040],seed[4029],seed[1154],seed[3403],seed[3593],seed[2972],seed[1297],seed[352],seed[2196],seed[1912],seed[2425],seed[2765],seed[3755],seed[1359],seed[1018],seed[359],seed[2204],seed[1735],seed[3927],seed[153],seed[787],seed[4048],seed[3748],seed[2517],seed[3164],seed[4068],seed[33],seed[3716],seed[4004],seed[2950],seed[795],seed[2708],seed[1344],seed[1443],seed[2267],seed[1317],seed[1070],seed[3267],seed[1533],seed[4028],seed[2615],seed[2370],seed[1095],seed[2392],seed[2036],seed[3817],seed[1522],seed[1930],seed[3498],seed[3934],seed[754],seed[2987],seed[2739],seed[642],seed[1838],seed[331],seed[2916],seed[1404],seed[518],seed[1933],seed[3029],seed[1349],seed[3401],seed[628],seed[680],seed[763],seed[1447],seed[3224],seed[1160],seed[2887],seed[2636],seed[3886],seed[1939],seed[469],seed[1545],seed[3890],seed[3673],seed[1825],seed[4067],seed[2978],seed[1757],seed[1266],seed[2527],seed[344],seed[2158],seed[136],seed[917],seed[78],seed[403],seed[2178],seed[408],seed[2882],seed[10],seed[2354],seed[2086],seed[3873],seed[69],seed[529],seed[701],seed[208],seed[3501],seed[34],seed[2531],seed[2287],seed[3249],seed[1026],seed[3888],seed[789],seed[792],seed[2157],seed[4018],seed[2378],seed[1798],seed[633],seed[2457],seed[2500],seed[3278],seed[435],seed[793],seed[1459],seed[526],seed[2989],seed[525],seed[209],seed[3588],seed[3907],seed[851],seed[429],seed[1902],seed[3519],seed[1102],seed[1839],seed[908],seed[2889],seed[1604],seed[1186],seed[3032],seed[2886],seed[2075],seed[3333],seed[107],seed[188],seed[1881],seed[1595],seed[324],seed[3713],seed[1040],seed[618],seed[886],seed[575],seed[211],seed[131],seed[2081],seed[3416],seed[3536],seed[67],seed[993],seed[961],seed[3611],seed[3814],seed[2830],seed[530],seed[196],seed[3766],seed[1988],seed[2728],seed[2984],seed[3859],seed[1059],seed[3439],seed[3304],seed[531],seed[1906],seed[2798],seed[1674],seed[2908],seed[3145],seed[678],seed[2911],seed[1634],seed[3273],seed[1851],seed[681],seed[1446],seed[3417],seed[2736],seed[3374],seed[2439],seed[3500],seed[1239],seed[466],seed[1201],seed[742],seed[1471],seed[2228],seed[629],seed[1190],seed[3894],seed[1931],seed[957],seed[2121],seed[1559],seed[645],seed[3446],seed[1363],seed[3453],seed[1943],seed[2324],seed[968],seed[1233],seed[1613],seed[3470],seed[2520],seed[3138],seed[3496],seed[1525],seed[3599],seed[747],seed[1206],seed[288],seed[256],seed[3441],seed[1509],seed[140],seed[1249],seed[2014],seed[2847],seed[2623],seed[1304],seed[520],seed[3572],seed[3734],seed[1842],seed[2330],seed[2526],seed[1341],seed[1272],seed[3187],seed[2415],seed[2738],seed[230],seed[1395],seed[1987],seed[3041],seed[467],seed[684],seed[105],seed[12],seed[3158],seed[303],seed[1913],seed[294],seed[3595],seed[3580],seed[3],seed[951],seed[3574],seed[2575],seed[1243],seed[1486],seed[1834],seed[3003],seed[2275],seed[2091],seed[816],seed[14],seed[339],seed[1847],seed[2203],seed[1647],seed[2676],seed[3113],seed[523],seed[1397],seed[3798],seed[2729],seed[2602],seed[2923],seed[3913],seed[1985],seed[1563],seed[2408],seed[4001],seed[1492],seed[941],seed[1106],seed[190],seed[4033],seed[1130],seed[1547],seed[551],seed[277],seed[1889],seed[2338],seed[2667],seed[900],seed[1997],seed[219],seed[312],seed[1136],seed[3456],seed[1739],seed[2928],seed[427],seed[1966],seed[2332],seed[267],seed[603],seed[2379],seed[167],seed[594],seed[1150],seed[3343],seed[519],seed[1683],seed[1978],seed[2760],seed[2162],seed[2404],seed[2762],seed[2835],seed[1333],seed[280],seed[2029],seed[3575],seed[1510],seed[953],seed[4088],seed[2302],seed[438],seed[4065],seed[2771],seed[1950],seed[343],seed[2349],seed[3603],seed[712],seed[3989],seed[1762],seed[1032],seed[18],seed[977],seed[1483],seed[3420],seed[3924],seed[315],seed[3825],seed[2595],seed[1846],seed[2910],seed[301],seed[1741],seed[2512],seed[2455],seed[859],seed[1806],seed[3657],seed[1539],seed[895],seed[2295],seed[2319],seed[2783],seed[1594],seed[3265],seed[1320],seed[3773],seed[3302],seed[3597],seed[3645],seed[1526],seed[2694],seed[2185],seed[1074],seed[4011],seed[1843],seed[2306],seed[989],seed[2871],seed[2627],seed[1809],seed[3505],seed[2549],seed[685],seed[599],seed[2990],seed[973],seed[2852],seed[95],seed[3561],seed[2460],seed[3976],seed[173],seed[36],seed[1515],seed[1265],seed[370],seed[2732],seed[2219],seed[812],seed[2447],seed[597],seed[2312],seed[260],seed[2441],seed[1161],seed[1462],seed[2993],seed[627],seed[3303],seed[814],seed[1294],seed[1875],seed[3843],seed[1714],seed[1772],seed[3436],seed[434],seed[1529],seed[3445],seed[4003],seed[2135],seed[3694],seed[1876],seed[2484],seed[2027],seed[2296],seed[1151],seed[2700],seed[753],seed[16],seed[3757],seed[2860],seed[1873],seed[2599],seed[1008],seed[1401],seed[3162],seed[1558],seed[2045],seed[1168],seed[2122],seed[975],seed[3393],seed[829],seed[1569],seed[2340],seed[3877],seed[616],seed[3384],seed[515],seed[2276],seed[3076],seed[1478],seed[4053],seed[1561],seed[1436],seed[2400],seed[3370],seed[1377],seed[2658],seed[2125],seed[1700],seed[2797],seed[3534],seed[317],seed[1699],seed[3607],seed[1895],seed[3939],seed[1188],seed[2977],seed[1226],seed[892],seed[3805],seed[316],seed[841],seed[871],seed[120],seed[2107],seed[3804],seed[2968],seed[746],seed[1274],seed[562],seed[117],seed[2854],seed[1348],seed[1612],seed[266],seed[868],seed[3360],seed[1835],seed[2969],seed[415],seed[2335],seed[547],seed[2689],seed[929],seed[3231],seed[1915],seed[3975],seed[2069],seed[1468],seed[456],seed[1830],seed[2813],seed[3533],seed[1463],seed[3233],seed[25],seed[1223],seed[440],seed[728],seed[411],seed[3788],seed[3553],seed[1244],seed[1474],seed[3083],seed[3627],seed[2453],seed[3925],seed[3021],seed[2022],seed[943],seed[985],seed[2190],seed[2872],seed[1788],seed[2795],seed[561],seed[827],seed[2681],seed[3022],seed[3062],seed[463],seed[3560],seed[1543],seed[302],seed[1110],seed[2628],seed[253],seed[1606],seed[1598],seed[1291],seed[788],seed[3653],seed[103],seed[4056],seed[3316],seed[3524],seed[3214],seed[2937],seed[2384],seed[306],seed[2181],seed[2412],seed[528],seed[3452],seed[43],seed[3831],seed[1019],seed[3151],seed[2539],seed[3306],seed[1442],seed[2072],seed[308],seed[2361],seed[44],seed[1626],seed[1068],seed[3232],seed[2980],seed[2294],seed[1221],seed[1975],seed[3320],seed[1012],seed[815],seed[3090],seed[1910],seed[2470],seed[579],seed[1343],seed[3209],seed[919],seed[1437],seed[3291],seed[1425],seed[174],seed[1952],seed[2868],seed[830],seed[2901],seed[3661],seed[590],seed[3218],seed[222],seed[3863],seed[2469],seed[2272],seed[735],seed[220],seed[2202],seed[3849],seed[3717],seed[2226],seed[1925],seed[3997],seed[1083],seed[1645],seed[675],seed[283],seed[844],seed[1681],seed[1819],seed[1938],seed[3827],seed[2982],seed[2318],seed[202],seed[3153],seed[2194],seed[2345],seed[273],seed[4015],seed[3821],seed[3747],seed[1560],seed[2610],seed[3590],seed[2925],seed[35],seed[3967],seed[1833],seed[233],seed[3811],seed[2479],seed[265],seed[803],seed[412],seed[3577],seed[1702],seed[1665],seed[2503],seed[444],seed[3922],seed[544],seed[2921],seed[905],seed[2633],seed[1776],seed[3485],seed[1310],seed[2971],seed[883],seed[1789],seed[4002],seed[2711],seed[2853],seed[175],seed[394],seed[1067],seed[2747],seed[1815],seed[1386],seed[3053],seed[3951],seed[171],seed[3292],seed[3495],seed[2101],seed[2104],seed[2954],seed[1078],seed[2433],seed[2616],seed[2806],seed[1305],seed[3228],seed[2651],seed[2594],seed[2822],seed[834],seed[620],seed[1995],seed[58],seed[2951],seed[1046],seed[1637],seed[1254],seed[1980],seed[3484],seed[1045],seed[1517],seed[39],seed[1077],seed[2848],seed[3276],seed[2037],seed[3486],seed[3672],seed[791],seed[2334],seed[181],seed[571],seed[3832],seed[1087],seed[1339],seed[1450],seed[3298],seed[3330],seed[3348],seed[1750],seed[2071],seed[3740],seed[1629],seed[672],seed[3902],seed[376],seed[1175],seed[3527],seed[655],seed[3957],seed[2932],seed[3014],seed[2170],seed[1361],seed[3425],seed[2111],seed[4066],seed[1063],seed[3647],seed[2067],seed[473],seed[4076],seed[799],seed[2857],seed[2252],seed[880],seed[1373],seed[3619],seed[3737],seed[2123],seed[3867],seed[3085],seed[221],seed[454],seed[2614],seed[102],seed[3404],seed[3891],seed[2592],seed[59],seed[566],seed[1421],seed[2945],seed[1648],seed[1234],seed[694],seed[3917],seed[1935],seed[1787],seed[2380],seed[3492],seed[4075],seed[311],seed[1718],seed[749],seed[45],seed[659],seed[2264],seed[3338],seed[2438],seed[138],seed[1156],seed[906],seed[1671],seed[3400],seed[2652],seed[2047],seed[364],seed[3082],seed[1192],seed[2829],seed[609],seed[619],seed[3736],seed[4077],seed[3389],seed[925],seed[1897],seed[1155],seed[3963],seed[739],seed[2746],seed[3034],seed[3613],seed[3691],seed[1752],seed[2348],seed[1023],seed[1942],seed[1917],seed[1860],seed[291],seed[2544],seed[564],seed[1241],seed[3714],seed[1643],seed[1736],seed[2501],seed[362],seed[3440],seed[205],seed[3379],seed[3764],seed[4034],seed[3852],seed[240],seed[3216],seed[3974],seed[3487],seed[3129],seed[481],seed[499],seed[3668],seed[3410],seed[305],seed[2618],seed[3357],seed[3217],seed[1774],seed[422],seed[1587],seed[1524],seed[313],seed[4085],seed[3636],seed[605],seed[1608],seed[1928],seed[1189],seed[2054],seed[3336],seed[3067],seed[1962],seed[1108],seed[1289],seed[3020],seed[3068],seed[2714],seed[1124],seed[2401],seed[3006],seed[3469],seed[3756],seed[2986],seed[4078],seed[1231],seed[2817],seed[1103],seed[1113],seed[607],seed[1396],seed[1368],seed[1242],seed[3666],seed[2118],seed[2748],seed[2959],seed[1213],seed[248],seed[3376],seed[3637],seed[3937],seed[3301],seed[4061],seed[166],seed[84],seed[3868],seed[1292],seed[3632],seed[3526],seed[580],seed[3172],seed[1378],seed[3133],seed[3194],seed[1552],seed[634],seed[955],seed[1687],seed[3464],seed[75],seed[2326],seed[121],seed[1281],seed[1355],seed[1017],seed[2686],seed[281],seed[3841],seed[836],seed[650],seed[2961],seed[1677],seed[3882],seed[1022],seed[2193],seed[2492],seed[432],seed[2612],seed[3378],seed[477],seed[2286],seed[3514],seed[1749],seed[660],seed[904],seed[3508],seed[3258],seed[2754],seed[2119],seed[262],seed[549],seed[3516],seed[1753],seed[3792],seed[3898],seed[3284],seed[326],seed[2182],seed[193],seed[360],seed[3846],seed[1465],seed[3406],seed[4019],seed[2692],seed[296],seed[2825],seed[1069],seed[805],seed[2581],seed[1163],seed[2973],seed[1907],seed[3328],seed[1250],seed[1432],seed[3537],seed[764],seed[1285],seed[1248],seed[3933],seed[2148],seed[2743],seed[237],seed[249],seed[1998],seed[1590],seed[1400],seed[3916],seed[2828],seed[1573],seed[2270],seed[1863],seed[3098],seed[1205],seed[3550],seed[2884],seed[322],seed[3540],seed[1521],seed[1593],seed[1801],seed[346],seed[48],seed[3159],seed[1454],seed[2976],seed[2502],seed[2198],seed[3725],seed[82],seed[1481],seed[7],seed[2629],seed[3033],seed[2019],seed[1507],seed[3184],seed[1885],seed[3354],seed[503],seed[2314],seed[3528],seed[1794],seed[3625],seed[4069],seed[3230],seed[3656],seed[704],seed[2533],seed[2476],seed[1399],seed[582],seed[1921],seed[3012],seed[976],seed[2768],seed[1831],seed[546],seed[3116],seed[4],seed[2468],seed[2056],seed[3325],seed[2095],seed[2154],seed[2396],seed[318],seed[270],seed[1007],seed[2559],seed[2924],seed[2706],seed[1477],seed[2998],seed[1945],seed[3010],seed[3066],seed[129],seed[2862],seed[3305],seed[722],seed[1423],seed[3319],seed[1879],seed[2292],seed[2547],seed[3142],seed[1968],seed[2508],seed[1754],seed[1607],seed[3879],seed[864],seed[1009],seed[2073],seed[417],seed[1636],seed[154],seed[2405],seed[2360],seed[3086],seed[2442],seed[3834],seed[2523],seed[1578],seed[148],seed[1107],seed[4047],seed[2756],seed[1491],seed[2558],seed[3810],seed[3568],seed[2981],seed[1790],seed[2970],seed[2366],seed[3576],seed[3799],seed[3893],seed[3600],seed[3803],seed[1245],seed[1461],seed[1005],seed[3418],seed[1054],seed[1194],seed[563],seed[765],seed[2192],seed[926],seed[2289],seed[1307],seed[1302],seed[3125],seed[289],seed[2929],seed[858],seed[3765],seed[3781],seed[806],seed[1235],seed[1695],seed[3490],seed[3398],seed[446],seed[1567],seed[1742],seed[1415],seed[299],seed[1716],seed[264],seed[538],seed[3875],seed[2514],seed[2015],seed[800],seed[3009],seed[3165],seed[1667],seed[2719],seed[2063],seed[398],seed[1411],seed[119],seed[4093],seed[2906],seed[2000],seed[3119],seed[643],seed[2661],seed[459],seed[1673],seed[3683],seed[1021],seed[3903],seed[1316],seed[3381],seed[527],seed[769],seed[2740],seed[3494],seed[1779],seed[2288],seed[1229],seed[2266],seed[995],seed[853],seed[1439],seed[3286],seed[4080],seed[3368],seed[334],seed[2807],seed[767],seed[3355],seed[77],seed[461],seed[949],seed[1963],seed[3429],seed[2551],seed[1941],seed[3155],seed[1125],seed[3178],seed[3107],seed[1455],seed[3570],seed[2861],seed[3995],seed[1610],seed[2042],seed[115],seed[2465],seed[179],seed[1803],seed[2787],seed[2565],seed[1094],seed[702],seed[2753],seed[3592],seed[287],seed[3851],seed[1694],seed[2087],seed[877],seed[1799],seed[3382],seed[1976],seed[3002],seed[258],seed[3708],seed[3272],seed[637],seed[2471],seed[3124],seed[1730],seed[2635],seed[3036],seed[513],seed[1661],seed[3684],seed[1375],seed[3709],seed[3587],seed[2168],seed[1185],seed[180],seed[197],seed[912],seed[76],seed[2299],seed[9],seed[683],seed[3136],seed[1015],seed[2698],seed[2483],seed[3615],seed[2026],seed[184],seed[1867],seed[1940],seed[2004],seed[132],seed[2274],seed[2053],seed[2572],seed[979],seed[1419],seed[843],seed[1624],seed[511],seed[3724],seed[68],seed[1269],seed[2995],seed[2790],seed[4009],seed[2939],seed[3548],seed[2632],seed[3941],seed[3222],seed[1965],seed[2333],seed[510],seed[176],seed[92],seed[2567],seed[4090],seed[3174],seed[711],seed[761],seed[768],seed[692],seed[3830],seed[2153],seed[2744],seed[474],seed[3866],seed[1715],seed[1565],seed[1562],seed[656],seed[1360],seed[2363],seed[1937],seed[3177],seed[888],seed[3435],seed[2530],seed[1807],seed[2391],seed[697],seed[654],seed[1982],seed[1322],seed[441],seed[165],seed[3839],seed[3602],seed[522],seed[653],seed[1713],seed[239],seed[2690],seed[1118],seed[1179],seed[2487],seed[1773],seed[1035],seed[2838],seed[4014],seed[991],seed[2061],seed[3881],seed[3118],seed[297],seed[885],seed[2488],seed[3651],seed[1719],seed[567],seed[2329],seed[1145],seed[1299],seed[2420],seed[2842],seed[472],seed[3442],seed[3763],seed[3361],seed[1109],seed[2562],seed[2003],seed[2017],seed[1449],seed[2328],seed[4021],seed[1698],seed[49],seed[2963],seed[1232],seed[3426],seed[2846],seed[3000],seed[1309],seed[191],seed[2824],seed[2648],seed[1866],seed[2207],seed[15],seed[1219],seed[2074],seed[2474],seed[1398],seed[228],seed[3309],seed[1336],seed[2452],seed[3397],seed[2879],seed[3812],seed[465],seed[1708],seed[3198],seed[416],seed[809],seed[61],seed[2209],seed[3658],seed[3678],seed[2702],seed[4007],seed[439],seed[3721],seed[2892],seed[1001],seed[2705],seed[1255],seed[2169],seed[2826],seed[2933],seed[3115],seed[1057],seed[1527],seed[2603],seed[1528],seed[2585],seed[2175],seed[1961],seed[1476],seed[101],seed[682],seed[3945],seed[2365],seed[2241],seed[2215],seed[3930],seed[1345],seed[2542],seed[2043],seed[504],seed[1922],seed[1193],seed[242],seed[1253],seed[1133],seed[1207],seed[341],seed[1936],seed[491],seed[507],seed[2305],seed[55],seed[1506],seed[4062],seed[3662],seed[3395],seed[3538],seed[1577],seed[1680],seed[4052],seed[1237],seed[2390],seed[2949],seed[1850],seed[2261],seed[897],seed[3789],seed[2406],seed[2269],seed[665],seed[971],seed[2774],seed[731],seed[1457],seed[2917],seed[996],seed[3451],seed[244],seed[2186],seed[2258],seed[1409],seed[1166],seed[948],seed[2358],seed[2236],seed[4020],seed[3955],seed[804],seed[2755],seed[4089],seed[201],seed[63],seed[2039],seed[3046],seed[1271],seed[719],seed[1775],seed[727],seed[2357],seed[3275],seed[1814],seed[862],seed[2089],seed[3065],seed[89],seed[3915],seed[1615],seed[2013],seed[1923],seed[2084],seed[218],seed[79],seed[1024],seed[2173],seed[2537],seed[3530],seed[3705],seed[4037],seed[486],seed[251],seed[23],seed[3205],seed[338],seed[2271],seed[3847],seed[2541],seed[676],seed[1746],seed[2229],seed[2115],seed[1918],seed[899],seed[2600],seed[3689],seed[1689],seed[3883],seed[1972],seed[2163],seed[3515],seed[480],seed[3001],seed[1920],seed[1117],seed[2232],seed[2254],seed[1004],seed[2426],seed[425],seed[389],seed[3711],seed[2735],seed[2421],seed[1508],seed[1066],seed[500],seed[3983],seed[4058],seed[570],seed[3506],seed[3285],seed[2934],seed[710],seed[3947],seed[3111],seed[2262],seed[3399],seed[73],seed[1887],seed[421],seed[3473],seed[3220],seed[268],seed[1261],seed[1137],seed[1721],seed[37],seed[2776],seed[3394],seed[3200],seed[2142],seed[1282],seed[2703],seed[667],seed[1784],seed[1592],seed[640],seed[3642],seed[3956],seed[3345],seed[720],seed[535],seed[3385],seed[2102],seed[1167],seed[1260],seed[3687],seed[1357],seed[3137],seed[2513],seed[3087],seed[2227],seed[2823],seed[2372],seed[2896],seed[1048],seed[3777],seed[3208],seed[4060],seed[790],seed[453],seed[3234],seed[1433],seed[766],seed[2076],seed[3535],seed[569],seed[3785],seed[688],seed[1640],seed[624],seed[3551],seed[1218],seed[1365],seed[1385],seed[3589],seed[3189],seed[3186],seed[1300],seed[3620],seed[20],seed[108],seed[2709],seed[2088],seed[122],seed[855],seed[125],seed[319],seed[2880],seed[1556],seed[3874],seed[2172],seed[4043],seed[447],seed[3547],seed[2282],seed[1127],seed[1581],seed[2213],seed[261],seed[2238],seed[2034],seed[658],seed[1816],seed[3655],seed[21],seed[1173],seed[2691],seed[2230],seed[541],seed[3402],seed[1099],seed[3288],seed[2516],seed[162],seed[1128],seed[3102],seed[212],seed[1381],seed[3173],seed[2371],seed[3612],seed[1489],seed[1389],seed[1583],seed[2991],seed[3202],seed[327],seed[884],seed[686],seed[2322],seed[357],seed[2831],seed[1039],seed[1430],seed[962],seed[1435],seed[3149],seed[3013],seed[1828],seed[3987],seed[3421],seed[3408],seed[3761],seed[3074],seed[3023],seed[3018],seed[3059],seed[3168],seed[568],seed[3140],seed[3801],seed[3112],seed[284],seed[1200],seed[2078],seed[2475],seed[2802],seed[88],seed[3984],seed[3105],seed[875],seed[1505],seed[3778],seed[785],seed[2313],seed[3386],seed[817],seed[2693],seed[2555],seed[1276],seed[2704],seed[4006],seed[1745],seed[243],seed[385],seed[2873],seed[810],seed[771],seed[2742],seed[966],seed[1956],seed[345],seed[3431],seed[2816],seed[2461],seed[1584],seed[3364],seed[1258],seed[1717],seed[3730],seed[1362],seed[1970],seed[1392],seed[198],seed[2440],seed[2489],seed[1871],seed[3281],seed[3324],seed[1536],seed[3921],seed[3938],seed[3206],seed[2291],seed[231],seed[3745],seed[3635],seed[178],seed[3121],seed[1198],seed[2504],seed[4071],seed[3608],seed[2145],seed[2553],seed[1888],seed[1662],seed[652],seed[1523],seed[1177],seed[3905],seed[4045],seed[104],seed[3850],seed[2161],seed[2875],seed[2779],seed[3936],seed[1599],seed[798],seed[2659],seed[661],seed[2660],seed[3719],seed[2930],seed[1537],seed[1981],seed[3299],seed[670],seed[2611],seed[2344],seed[1532],seed[2409],seed[2395],seed[2410],seed[350],seed[3567],seed[714],seed[3546],seed[707],seed[3466],seed[151],seed[2671],seed[2878],seed[410],seed[1143],seed[3317],seed[3741],seed[3271],seed[560],seed[1171],seed[1551],seed[2138],seed[3920],seed[2786],seed[65],seed[915],seed[826],seed[2552],seed[577],seed[3024],seed[2281],seed[3160],seed[2699],seed[2893],seed[1554],seed[3161],seed[3212],seed[247],seed[2350],seed[1418],seed[1056],seed[1600],seed[3563],seed[1726],seed[1657],seed[4079],seed[146],seed[2573],seed[2362],seed[3504],seed[2683],seed[3242],seed[2864],seed[1826],seed[3480],seed[2808],seed[3775],seed[1488],seed[3605],seed[2310],seed[3864],seed[3092],seed[3123],seed[870],seed[3353],seed[133],seed[2066],seed[2718],seed[748],seed[2948],seed[876],seed[1482],seed[1326],seed[3327],seed[337],seed[3463],seed[3910],seed[2979],seed[3918],seed[2710],seed[802],seed[2890],seed[3007],seed[1484],seed[657],seed[1652],seed[1518],seed[1631],seed[1856],seed[3562],seed[1511],seed[3372],seed[3210],seed[3630],seed[1767],seed[517],seed[3039],seed[1184],seed[646],seed[3641],seed[2940],seed[2863],seed[381],seed[1743],seed[130],seed[1142],seed[2277],seed[1350],seed[600],seed[1855],seed[46],seed[1055],seed[1804],seed[1479],seed[1911],seed[4040],seed[584],seed[255],seed[916],seed[3071],seed[689],seed[2459],seed[2195],seed[1722],seed[860],seed[782],seed[832],seed[1705],seed[3122],seed[3377],seed[1660],seed[537],seed[1327],seed[3088],seed[3986],seed[3307],seed[2759],seed[1230],seed[1646],seed[2577],seed[1215],seed[3289],seed[4082],seed[2877],seed[1601],seed[913],seed[3970],seed[2525],seed[3681],seed[2339],seed[2785],seed[3806],seed[3784],seed[1338],seed[846],seed[4027],seed[3179],seed[2761],seed[141],seed[3460],seed[1164],seed[1520],seed[3196],seed[2435],seed[323],seed[293],seed[2952],seed[2048],seed[87],seed[881],seed[3323],seed[3581],seed[762],seed[3979],seed[206],seed[3089],seed[2206],seed[3552],seed[458],seed[2033],seed[60],seed[1306],seed[2701],seed[2805],seed[155],seed[3972],seed[2545],seed[1513],seed[3467],seed[1312],seed[2355],seed[3751],seed[2256],seed[1901],seed[3294],seed[2912],seed[210],seed[2352],seed[585],seed[4070],seed[1546],seed[3326],seed[3128],seed[1793],seed[2598],seed[1603],seed[2393],seed[2347],seed[1737],seed[698],seed[3855],seed[3359],seed[1549],seed[428],seed[161],seed[1820],seed[558],seed[1622],seed[673],seed[2568],seed[1678],seed[3601],seed[1979],seed[1394],seed[1003],seed[2766],seed[669],seed[2308],seed[1633],seed[1666],seed[2092],seed[2490],seed[2343],seed[110],seed[3465],seed[1217],seed[71],seed[2472],seed[252],seed[2985],seed[1380],seed[588],seed[3621],seed[4054],seed[2609],seed[553],seed[2665],seed[2251],seed[1574],seed[200],seed[1458],seed[3176],seed[1079],seed[4064],seed[2764],seed[820],seed[2670],seed[887],seed[1440],seed[2085],seed[2788],seed[3080],seed[2211],seed[3097],seed[2664],seed[3491],seed[1865],seed[1621],seed[2607],seed[177],seed[1273],seed[118],seed[1720],seed[3900],seed[2116],seed[62],seed[1944],seed[1672],seed[573],seed[3130],seed[3223],seed[2590],seed[2321],seed[758],seed[1356],seed[1905],seed[2259],seed[3110],seed[2099],seed[3848],seed[3791],seed[935],seed[1490],seed[2159],seed[1036],seed[1061],seed[409],seed[2283],seed[796],seed[4087],seed[3943],seed[1420],seed[3558],seed[1605],seed[2300],seed[3297],seed[2891],seed[2216],seed[2515],seed[2280],seed[965],seed[1174],seed[1501],seed[550],seed[921],seed[911],seed[540],seed[375],seed[2898],seed[2369],seed[215],seed[1924],seed[625],seed[3019],seed[3409],seed[2141],seed[928],seed[2597],seed[2535],seed[460],seed[1596],seed[988],seed[3075],seed[2035],seed[3016],seed[647],seed[3557],seed[2257],seed[4013],seed[2849],seed[3419],seed[1031],seed[1303],seed[1050],seed[149],seed[3371],seed[1119],seed[111],seed[74],seed[2151],seed[1530],seed[3135],seed[3633],seed[3070],seed[156],seed[2639],seed[2682],seed[1453],seed[2713],seed[1759],seed[4072],seed[232],seed[4074],seed[3606],seed[2336],seed[38],seed[752],seed[2579],seed[1144],seed[1251],seed[1126],seed[2093],seed[2625],seed[3352],seed[1264],seed[2165],seed[3422],seed[2947],seed[3758],seed[325],seed[2070],seed[3675],seed[3591],seed[4050],seed[2375],seed[2136],seed[2593],seed[778],seed[1367],seed[986],seed[1279],seed[1747],seed[97],seed[3772],seed[3424],seed[3964],seed[246],seed[2543],seed[2315],seed[3704],seed[2117],seed[1585],seed[54],seed[2325],seed[424],seed[2255],seed[920],seed[361],seed[2578],seed[207],seed[2249],seed[4049],seed[3703],seed[2001],seed[128],seed[1116],seed[2411],seed[145],seed[506],seed[1785],seed[2407],seed[3583],seed[3807],seed[356],seed[2217],seed[1782],seed[3388],seed[775],seed[26],seed[592],seed[1899],seed[2673],seed[1211],seed[2994],seed[2874],seed[3996],seed[1731],seed[2399],seed[47],seed[304],seed[2902],seed[1542],seed[2707],seed[2630],seed[3434],seed[3503],seed[3197],seed[3030],seed[1620],seed[2131],seed[593],seed[3350],seed[1684],seed[3688],seed[992],seed[1602],seed[1131],seed[2587],seed[2750],seed[2794],seed[2678],seed[4035],seed[2905],seed[3497],seed[40],seed[3185],seed[2645],seed[1],seed[1157],seed[3259],seed[3433],seed[891],seed[2649],seed[3928],seed[3796],seed[3670],seed[2996],seed[565],seed[2058],seed[1777],seed[159],seed[2105],seed[3157],seed[2064],seed[1278],seed[777],seed[2278],seed[3269],seed[93],seed[2834],seed[2637],seed[937],seed[3407],seed[3489],seed[3525],seed[856],seed[2201],seed[2804],seed[1058],seed[2389],seed[3084],seed[534],seed[2051],seed[923],seed[2638],seed[2622],seed[1783],seed[1832],seed[1456],seed[2183],seed[1448],seed[1791],seed[1081],seed[3150],seed[548],seed[479],seed[2960],seed[1579],seed[1014],seed[351],seed[581],seed[1475],seed[1880],seed[3818],seed[4030],seed[1751],seed[476],seed[980],seed[3518],seed[1387],seed[1104],seed[2833],seed[1686],seed[1006],seed[3911],seed[3449],seed[1197],seed[332],seed[3493],seed[2810],seed[1796],seed[3573],seed[3985],seed[615],seed[1135],seed[2481],seed[2550],seed[3499],seed[743],seed[3366],seed[502],seed[2915],seed[1159],seed[1372],seed[1538],seed[418],seed[2049],seed[2723],seed[3582],seed[2443],seed[2770],seed[139],seed[2382],seed[2655],seed[2851],seed[85],seed[3935],seed[3586],seed[3152],seed[2999],seed[3896],seed[611],seed[2644],seed[3901],seed[2869],seed[2120],seed[2140],seed[1853],seed[2268],seed[3584],seed[613],seed[1960],seed[330],seed[1053],seed[42],seed[182],seed[1034],seed[1347],seed[2926],seed[2741],seed[505],seed[3646],seed[94],seed[2147],seed[773],seed[1216],seed[2446],seed[3697],seed[1894],seed[2096],seed[2936],seed[2643],seed[716],seed[137],seed[982],seed[2867],seed[2414],seed[865],seed[377],seed[2046],seed[328],seed[572],seed[1366],seed[3108],seed[1861],seed[1335],seed[2265],seed[2646],seed[2956],seed[533],seed[3191],seed[1374],seed[1948],seed[3731],seed[285],seed[1246],seed[3256],seed[2663],seed[3578],seed[1971],seed[750],seed[2006],seed[3254],seed[164],seed[436],seed[1844],seed[3332],seed[1916],seed[784],seed[3120],seed[1331],seed[397],seed[898],seed[3396],seed[852],seed[2495],seed[172],seed[371],seed[3968],seed[2941],seed[2028],seed[1065],seed[2641],seed[3695],seed[1572],seed[1890],seed[29],seed[170],seed[622],seed[1644],seed[954],seed[2528],seed[1120],seed[1692],seed[1874],seed[2221],seed[2858],seed[3529],seed[1813],seed[1738],seed[4055],seed[2773],seed[3203],seed[833],seed[934],seed[4023],seed[770],seed[1780],seed[2675],seed[612],seed[2604],seed[158],seed[1909],seed[1649],seed[3767],seed[759],seed[2983],seed[2243],seed[1575],seed[1016],seed[854],seed[3038],seed[751],seed[2927],seed[1727],seed[3669],seed[999],seed[2584],seed[3311],seed[3991],seed[217],seed[114],seed[3835],seed[3842],seed[3117],seed[1829],seed[2922],seed[3759],seed[1707],seed[873],seed[2463],seed[1115],seed[1139],seed[2818],seed[1550],seed[3443],seed[3824],seed[2456],seed[1852],seed[4084],seed[3474],seed[4008],seed[1140],seed[1002],seed[3664],seed[1709],seed[1823],seed[890],seed[946],seed[649],seed[2497],seed[124],seed[2129],seed[3415],seed[1351],seed[1632],seed[1228],seed[2137],seed[3049],seed[3942],seed[1369],seed[402],seed[3427],seed[2582],seed[3723],seed[390],seed[223],seed[1630],seed[3069],seed[3461],seed[1122],seed[3251],seed[3944],seed[2174],seed[2510],seed[1926],seed[369],seed[443],seed[3701],seed[2606],seed[2245],seed[2155],seed[3769],seed[1953],seed[2478],seed[3237],seed[863],seed[1358],seed[2052],seed[3280],seed[3965],seed[1676],seed[717],seed[2021],seed[3571],seed[1869],seed[3329],seed[2381],seed[1744],seed[3008],seed[1098],seed[3126],seed[942],seed[2684],seed[3405],seed[3509],seed[406],seed[1992],seed[559],seed[2397],seed[478],seed[3904],seed[1540],seed[2285],seed[163],seed[3783],seed[774],seed[3978],seed[1494],seed[1771],seed[2486],seed[3260],seed[3960],seed[157],seed[1900],seed[3005],seed[2975],seed[423],seed[970],seed[1121],seed[1332],seed[358],seed[3829],seed[3502],seed[1170],seed[744],seed[3610],seed[2509],seed[849],seed[2128],seed[857],seed[83],seed[981],seed[664],seed[1041],seed[1723],seed[1974],seed[320],seed[1202],seed[2812],seed[578],seed[471],seed[3238],seed[3629],seed[2246],seed[1408],seed[3423],seed[932],seed[2342],seed[2965],seed[1765],seed[1576],seed[3981],seed[1262],seed[1841],seed[1199],seed[963],seed[2388],seed[1178],seed[2666],seed[2796],seed[2210],seed[1247],seed[3457],seed[1623],seed[3523],seed[3786],seed[3127],seed[772],seed[691],seed[2799],seed[2466],seed[3828],seed[1405],seed[1802],seed[395],seed[99],seed[690],seed[2712],seed[2653],seed[2367],seed[455],seed[1589],seed[1864],seed[958],seed[2149],seed[1642],seed[1499],seed[997],seed[3585],seed[3390],seed[1996],seed[3143],seed[2913],seed[4017],seed[3148],seed[2844],seed[1792],seed[3363],seed[1183],seed[2467],seed[194],seed[2214],seed[3753],seed[3845],seed[1428],seed[3468],seed[1180],seed[1010],seed[3926],seed[1821],seed[2674],seed[70],seed[3109],seed[2942],seed[1653],seed[3296],seed[626],seed[1770],seed[1298],seed[2260],seed[1973],seed[2044],seed[3091],seed[726],seed[1984],seed[1187],seed[2687],seed[2177],seed[2018],seed[2726],seed[2730],seed[2082],seed[3543],seed[2250],seed[1346],seed[309],seed[238],seed[2364],seed[3762],seed[2445],seed[1704],seed[3887],seed[894],seed[493],seed[3980],seed[1132],seed[3351],seed[1516],seed[2432],seed[4092],seed[2914],seed[3063],seed[3510],seed[1641],seed[374],seed[909],seed[143],seed[2077],seed[2885],seed[2020],seed[3660],seed[3726],seed[3282],seed[824],seed[2919],seed[1256],seed[3954],seed[2057],seed[2524],seed[28],seed[3609],seed[1325],seed[2002],seed[3884],seed[1487],seed[1854],seed[3895],seed[2112],seed[2784],seed[2431],seed[1496],seed[2668],seed[3802],seed[2007],seed[1849],seed[2040],seed[2506],seed[1123],seed[3146],seed[524],seed[2309],seed[1165],seed[1733],seed[757],seed[51],seed[2132],seed[2290],seed[80],seed[3952],seed[604],seed[952],seed[3872],seed[2114],seed[3973],seed[3414],seed[1000],seed[3545],seed[2180],seed[866],seed[3513],seed[536],seed[3225],seed[1480],seed[3702],seed[3483],seed[1434],seed[552],seed[4036],seed[1227],seed[4073],seed[1568],seed[3686],seed[1729],seed[2647],seed[213],seed[3556],seed[462],seed[2688],seed[1275],seed[1701],seed[556],seed[2143],seed[3696],seed[383],seed[3077],seed[2957],seed[3204],seed[677],seed[1426],seed[606],seed[8],seed[848],seed[4005],seed[1402],seed[1416],seed[2560],seed[1208],seed[614],seed[3857],seed[32],seed[2331],seed[1314],seed[1321],seed[1580],seed[3195],seed[2403],seed[3247],seed[3682],seed[274],seed[4086],seed[3035],seed[674],seed[3060],seed[401],seed[3261],seed[1500],seed[2962],seed[2621],seed[1444],seed[1495],seed[3101],seed[2782],seed[1582],seed[3690],seed[1502],seed[3383],seed[407],seed[1711],seed[1076],seed[2303],seed[709],seed[3707],seed[98],seed[127],seed[382],seed[1553],seed[1761],seed[2394],seed[2809],seed[5],seed[3134],seed[2566],seed[3347],seed[2832],seed[2197],seed[3450],seed[3746],seed[1818],seed[3680],seed[2840],seed[1284],seed[1836],seed[3643],seed[2450],seed[1725],seed[1519],seed[3293],seed[2424],seed[708],seed[984],seed[1288],seed[1364],seed[3058],seed[3950],seed[1101],seed[354],seed[1685],seed[3335],seed[2376],seed[189],seed[3892],seed[22],seed[3880],seed[2184],seed[4057],seed[699],seed[2247],seed[3213],seed[497],seed[601],seed[922],seed[3430],seed[1295],seed[2897],seed[66],seed[1267],seed[3055],seed[2242],seed[3428],seed[1146],seed[109],seed[1617],seed[2298],seed[286],seed[3050],seed[1152],seed[1668],seed[1859],seed[336],seed[2098],seed[3479],seed[3663],seed[695],seed[2359],seed[3444],seed[2301],seed[1712],seed[1445],seed[451],seed[185],seed[718],seed[2751],seed[431],seed[3631],seed[3246],seed[3649],seed[1564],seed[1195],seed[3056],seed[896],seed[2423],seed[3215],seed[147],seed[91],seed[2297],seed[3840],seed[1503],seed[3899],seed[3932],seed[840],seed[2697],seed[2152],seed[426],seed[1393],seed[2430],seed[4010],seed[3257],seed[1635],seed[380],seed[31],seed[367],seed[2904],seed[3738],seed[780],seed[1379],seed[353],seed[1096],seed[3712],seed[3072],seed[187],seed[64],seed[1220],seed[2279],seed[3478],seed[3760],seed[2133],seed[2669],seed[1654],seed[1090],seed[2496],seed[783],seed[1703],seed[3106],seed[3644],seed[1959],seed[1340],seed[2589],seed[3315],seed[1371],seed[2617],seed[2224],seed[3774],seed[314],seed[776],seed[532],seed[276],seed[494],seed[3253],seed[2103],seed[241],seed[3241],seed[1138],seed[1786],seed[1293],seed[3201],seed[631],seed[250],seed[2888],seed[1105],seed[1656],seed[1033],seed[1758],seed[2819],seed[1388],seed[144],seed[740],seed[2856],seed[1958],seed[1071],seed[960],seed[2387],seed[2850],seed[3331],seed[1051],seed[3373],seed[2008],seed[2841],seed[365],seed[3517],seed[3750],seed[1679],seed[52],seed[1319],seed[399],seed[3797],seed[2437],seed[19],seed[1919],seed[457],seed[910],seed[967],seed[271],seed[2032],seed[2767],seed[1691],seed[1877],seed[482],seed[1964],seed[1311],seed[1999],seed[823],seed[2055],seed[4024],seed[1280],seed[2583],seed[2845],seed[555],seed[666],seed[3263],seed[86],seed[2814],seed[3219],seed[3511],seed[3953],seed[760],seed[610],seed[1993],seed[279],seed[3626],seed[414],seed[3624],seed[3961],seed[2449],seed[3476],seed[100],seed[3015],seed[468],seed[721],seed[2988],seed[1728],seed[2222],seed[737],seed[3349],seed[514],seed[3477],seed[1892],seed[2187],seed[1862],seed[3815],seed[0],seed[2576],seed[2791],seed[1891],seed[90],seed[2827],seed[1498],seed[4039],seed[168],seed[1591],seed[847],seed[3472],seed[2494],seed[930],seed[3833],seed[2758],seed[419],seed[2124],seed[630],seed[1286],seed[1983],seed[2716],seed[1619],seed[1296],seed[3539],seed[3794],seed[703],seed[3095],seed[2083],seed[2402],seed[1812],seed[1990],seed[2263],seed[1706],seed[1955],seed[1422],seed[3226],seed[2160],seed[501],seed[134],seed[321],seed[17],seed[3598],seed[1093],seed[3971],seed[387],seed[1270],seed[1535],seed[3982],seed[3365],seed[2239],seed[2997],seed[822],seed[496],seed[1967],seed[2024],seed[3969],seed[723],seed[907],seed[3648],seed[290],seed[2657],seed[2068],seed[3268],seed[4044],seed[263],seed[1756],seed[745],seed[1473],seed[2538],seed[1566],seed[2591],seed[2200],seed[1470],seed[1655],seed[2775],seed[275],seed[3236],seed[413],seed[2859],seed[490],seed[2094],seed[3054],seed[126],seed[442],seed[786],seed[1329],seed[1224],seed[2554],seed[3240],seed[2640],seed[2821],seed[1072],seed[1181],seed[1886],seed[819],seed[1466],seed[2752],seed[1534],seed[3958],seed[2564],seed[2870],seed[57],seed[3674],seed[2757],seed[2059],seed[3166],seed[4032],seed[214],seed[869],seed[1318],seed[861],seed[2171],seed[2866],seed[781],seed[587],seed[1932],seed[1469],seed[940],seed[292],seed[2521],seed[3369],seed[730],seed[1618],seed[498],seed[3042],seed[3531],seed[1337],seed[2793],seed[282],seed[3132],seed[3507],seed[2626],seed[3052],seed[2451],seed[1027],seed[3808],seed[4012],seed[3940],seed[1734],seed[2580],seed[3617],seed[3180],seed[386],seed[1313],seed[4083],seed[2134],seed[342],seed[3715],seed[1805],seed[388],seed[470],seed[192],seed[363],seed[3448],seed[1080],seed[1342],seed[1732],seed[2100],seed[234],seed[1969],seed[2769],seed[2248],seed[1088],seed[641],seed[2938],seed[3865],seed[1858],seed[1989],seed[1611],seed[3182],seed[2030],seed[1410],seed[1609],seed[3459],seed[1100],seed[2419],seed[1837],seed[1196],seed[1268],seed[3650],seed[2418],seed[671],seed[3768],seed[3838],seed[2571],seed[3047],seed[1659],seed[2188],seed[1638],seed[825],seed[3078],seed[1413],seed[2815],seed[3412],seed[1724],seed[2781],seed[450],seed[2493],seed[554],seed[2434],seed[2284],seed[3290],seed[1898],seed[1169],seed[1896],seed[2534],seed[3819],seed[3048],seed[379],seed[3754],seed[2144],seed[3885],seed[3156],seed[1162],seed[1760],seed[3638],seed[3011],seed[3685],seed[2462],seed[3114],seed[974],seed[340],seed[3057],seed[3856],seed[1020],seed[3262],seed[1062],seed[2353],seed[794],seed[2025],seed[1158],seed[3988],seed[1639],seed[2237],seed[1287],seed[2079],seed[226],seed[639],seed[2016],seed[3622],seed[3949],seed[1977],seed[1808],seed[3447],seed[4025],seed[1778],seed[2800],seed[2205],seed[1810],seed[3919],seed[1148],seed[2108],seed[1429],seed[2060],seed[2955],seed[2772],seed[1914],seed[1893],seed[3342],seed[3235],seed[3722],seed[2642],seed[1240],seed[1822],seed[245],seed[938],seed[994],seed[2212],seed[2920],seed[3618],seed[635],seed[1927],seed[713],seed[3340],seed[3853],seed[2304],seed[2398],seed[3163],seed[3028],seed[1710],seed[3521],seed[2199],seed[2065],seed[2307],seed[169],seed[3227],seed[3923],seed[1354],seed[3718],seed[3044],seed[1176],seed[4038],seed[1334],seed[2634],seed[464],seed[3889],seed[2724],seed[3099],seed[3244],seed[3728],seed[1878],seed[225],seed[1840],seed[3252],seed[596],seed[4031],seed[2820],seed[2803],seed[1212],seed[2620],seed[1857],seed[3094],seed[2233],seed[729],seed[310],seed[1441],seed[135],seed[487],seed[3471],seed[3239],seed[56],seed[4081],seed[348],seed[2253],seed[3813],seed[2903],seed[959],seed[3671],seed[1464],seed[2139],seed[874],seed[2416],seed[4042],seed[1570],seed[2778],seed[903],seed[6],seed[492],seed[1497],seed[2725],seed[914],seed[2749],seed[3387],seed[944],seed[2540],seed[333],seed[2931],seed[3634],seed[839],seed[1755],seed[2377],seed[1149],seed[2511],seed[186],seed[3579],seed[1616],seed[828],seed[3270],seed[3248],seed[638],seed[3541],seed[2320],seed[229],seed[195],seed[2966],seed[838],seed[4000],seed[3064],seed[3793],seed[235],seed[3188],seed[3732],seed[366],seed[3549],seed[2235],seed[3854],seed[50],seed[2429],seed[3481],seed[3512],seed[983],seed[2624],seed[483],seed[433],seed[2491],seed[1693],seed[437],seed[2146],seed[1817],seed[648],seed[3522],seed[3770],seed[3154],seed[4091],seed[2482],seed[3959],seed[3308],seed[1951],seed[508],seed[927],seed[700],seed[2715],seed[2127],seed[2876],seed[574],seed[2485],seed[632],seed[545],seed[3169],seed[3520],seed[893],seed[1669],seed[801],seed[485],seed[378],seed[2546],seed[1407],seed[668],seed[608],seed[3314],seed[495],seed[1204],seed[2386],seed[3998],seed[2680],seed[3131],seed[589],seed[3043],seed[1748],seed[3679],seed[3183],seed[1845],seed[2569],seed[3141],seed[3614],seed[2518],seed[889],seed[2507],seed[3604],seed[3344],seed[2413],seed[2522],seed[2570],seed[3897],seed[3809],seed[1089],seed[3749],seed[224],seed[3966],seed[808],seed[400],seed[3596],seed[3300],seed[368],seed[1904],seed[2351],seed[3826],seed[1827],seed[1903],seed[1403],seed[2935],seed[2992],seed[2631],seed[449],seed[1203],seed[1682],seed[2010],seed[2696],seed[3735],seed[2722],seed[2422],seed[998],seed[3594],seed[3729],seed[1236],seed[969],seed[1086],seed[4051],seed[3190],seed[1627],seed[842],seed[939],seed[3667],seed[2720],seed[850],seed[595],seed[2601],seed[3565],seed[1052],seed[872],seed[2505],seed[696],seed[3266],seed[705],seed[1028],seed[2041],seed[2519],seed[1571],seed[1994],seed[3167],seed[679],seed[2317],seed[4026],seed[2946],seed[2909],seed[2717],seed[3743],seed[3004],seed[3287],seed[1324],seed[3193],seed[598],seed[1047],seed[3475],seed[1848],seed[918],seed[724],seed[3367],seed[3455],seed[2189],seed[3488],seed[924],seed[2385],seed[1811],seed[2605],seed[183],seed[2792],seed[2974],seed[430],seed[2672],seed[1214],seed[3640],seed[583],seed[3836],seed[1084],seed[3569],seed[1222],seed[2130],seed[931],seed[1493],seed[3337],seed[2080],seed[272],seed[2900],seed[3909],seed[4095],seed[2374],seed[1868],seed[349],seed[204],seed[160],seed[2498],seed[2427],seed[3375],seed[3250],seed[257],seed[2839],seed[1555],seed[978],seed[3871],seed[355],seed[1182],seed[3931],seed[488],seed[3860],seed[1438],seed[1301],seed[557],seed[3665],seed[106],seed[1097],seed[1472],seed[807],seed[295],seed[254],seed[335],seed[3199],seed[2480],seed[2695],seed[445],seed[1797],seed[3380],seed[1658],seed[3221],seed[2327],seed[1384],seed[2323],seed[4094],seed[687],seed[3341],seed[3906],seed[259],seed[964],seed[1514],seed[3559],seed[2958],seed[1541],seed[2223],seed[2588],seed[3277],seed[693],seed[2685],seed[756],seed[3908],seed[818],seed[1044],seed[2731],seed[2106],seed[3139],seed[3554],seed[797],seed[3192],seed[4041],seed[1075],seed[835],seed[2737],seed[1986],seed[2031],seed[1414],seed[1544],seed[203],seed[2417],seed[3283],seed[3482],seed[1586],seed[3800],seed[3312],seed[1064],seed[1290],seed[3318],seed[663],seed[3073],seed[1690],seed[3771],seed[393],seed[3977],seed[2943],seed[3313],seed[779],seed[2536],seed[2150],seed[24],seed[3555],seed[404],seed[878],seed[4016],seed[3790],seed[2557],seed[2734],seed[1112],seed[3170],seed[405],seed[3795],seed[3623],seed[3566],seed[2477],seed[1025],seed[3310],seed[1697],seed[1370],seed[1073],seed[1460],seed[2341],seed[2464],seed[1884],seed[3844],seed[2473],seed[2368],seed[1947],seed[3742],seed[1049],seed[1315],seed[1085],seed[199],seed[516],seed[1650],seed[1504],seed[2881],seed[755],seed[3362],seed[3322],seed[1323],seed[586],seed[2244],seed[3438],seed[3659],seed[956],seed[2428],seed[269],seed[901],seed[3994],seed[1383],seed[2126],seed[3181],seed[1766],seed[3876],seed[3992],seed[1991],seed[3391],seed[2733],seed[1153],seed[1134],seed[2837],seed[2855],seed[2062],seed[152],seed[1946],seed[950],seed[448],seed[1424],seed[3948],seed[2780],seed[3229],seed[2899],seed[3744],seed[2918]}; 
//        seed6 <= {seed[3333],seed[1882],seed[2180],seed[1478],seed[347],seed[3824],seed[9],seed[1363],seed[1908],seed[2134],seed[2917],seed[2601],seed[4038],seed[2948],seed[3576],seed[2516],seed[3599],seed[1370],seed[1913],seed[1089],seed[3313],seed[1462],seed[2216],seed[492],seed[1912],seed[1024],seed[3045],seed[3510],seed[909],seed[252],seed[3377],seed[3179],seed[587],seed[1482],seed[1396],seed[1835],seed[1866],seed[1997],seed[1278],seed[2660],seed[2382],seed[851],seed[3964],seed[1839],seed[2447],seed[2776],seed[864],seed[3194],seed[680],seed[359],seed[613],seed[1410],seed[1124],seed[2529],seed[2806],seed[3679],seed[3043],seed[519],seed[2589],seed[2804],seed[4050],seed[1394],seed[1144],seed[161],seed[125],seed[767],seed[3307],seed[4082],seed[2977],seed[2003],seed[3253],seed[4077],seed[3471],seed[3230],seed[3488],seed[154],seed[2843],seed[3072],seed[1443],seed[3055],seed[1461],seed[1915],seed[1353],seed[1250],seed[1006],seed[2118],seed[3139],seed[2068],seed[1776],seed[1179],seed[4063],seed[3823],seed[1760],seed[972],seed[391],seed[2527],seed[726],seed[228],seed[112],seed[245],seed[500],seed[1115],seed[3845],seed[581],seed[1890],seed[2803],seed[429],seed[2832],seed[2787],seed[870],seed[3787],seed[3640],seed[3722],seed[2188],seed[461],seed[2793],seed[1301],seed[2288],seed[2189],seed[2570],seed[3171],seed[2822],seed[3478],seed[3835],seed[3792],seed[298],seed[3019],seed[3553],seed[2362],seed[50],seed[3669],seed[1509],seed[3033],seed[1737],seed[1031],seed[1649],seed[3305],seed[3991],seed[1495],seed[1650],seed[2119],seed[771],seed[2884],seed[2503],seed[2786],seed[617],seed[3858],seed[1824],seed[1429],seed[596],seed[996],seed[46],seed[1576],seed[232],seed[559],seed[85],seed[974],seed[3592],seed[1075],seed[2468],seed[1718],seed[3147],seed[3632],seed[1813],seed[3736],seed[1193],seed[4040],seed[3409],seed[3235],seed[1800],seed[2761],seed[676],seed[1874],seed[3187],seed[1052],seed[2092],seed[1037],seed[3495],seed[1397],seed[2359],seed[631],seed[2102],seed[643],seed[2878],seed[4011],seed[2038],seed[3695],seed[3862],seed[2401],seed[2831],seed[1766],seed[714],seed[3976],seed[1785],seed[355],seed[3001],seed[2421],seed[1816],seed[1349],seed[250],seed[1273],seed[2735],seed[3412],seed[1811],seed[3830],seed[2290],seed[1696],seed[1621],seed[964],seed[3343],seed[1023],seed[2056],seed[1610],seed[3786],seed[1085],seed[2898],seed[2683],seed[2959],seed[603],seed[1653],seed[2133],seed[2823],seed[799],seed[3838],seed[2517],seed[3465],seed[3366],seed[3295],seed[3829],seed[3500],seed[2053],seed[3827],seed[2173],seed[2954],seed[947],seed[3924],seed[3586],seed[2870],seed[2961],seed[1065],seed[2137],seed[418],seed[442],seed[128],seed[313],seed[1463],seed[898],seed[1294],seed[412],seed[2398],seed[991],seed[1266],seed[1688],seed[2992],seed[755],seed[3116],seed[258],seed[805],seed[3330],seed[2923],seed[2391],seed[3997],seed[3698],seed[3107],seed[1487],seed[163],seed[1257],seed[2183],seed[1859],seed[143],seed[3565],seed[139],seed[1377],seed[3548],seed[3590],seed[1526],seed[748],seed[2984],seed[3987],seed[3185],seed[1472],seed[3563],seed[3146],seed[259],seed[620],seed[4062],seed[1086],seed[2711],seed[1585],seed[957],seed[2349],seed[1909],seed[1947],seed[2813],seed[3387],seed[2494],seed[2629],seed[2333],seed[2368],seed[2895],seed[2700],seed[3371],seed[3690],seed[1562],seed[990],seed[1427],seed[3524],seed[1697],seed[281],seed[80],seed[2544],seed[1107],seed[2689],seed[4078],seed[529],seed[1473],seed[2669],seed[1035],seed[3110],seed[1453],seed[1715],seed[2746],seed[4047],seed[200],seed[2591],seed[155],seed[1063],seed[3952],seed[1387],seed[1214],seed[3340],seed[1860],seed[3096],seed[448],seed[4018],seed[1351],seed[1002],seed[3130],seed[2040],seed[4004],seed[2723],seed[3948],seed[1659],seed[286],seed[2587],seed[89],seed[60],seed[2267],seed[1008],seed[1259],seed[3250],seed[826],seed[2082],seed[850],seed[2900],seed[215],seed[253],seed[729],seed[1579],seed[3483],seed[1440],seed[3456],seed[761],seed[1428],seed[1941],seed[1522],seed[815],seed[2017],seed[1898],seed[1442],seed[2208],seed[2159],seed[3814],seed[1729],seed[3803],seed[3405],seed[892],seed[396],seed[1983],seed[1437],seed[3419],seed[3125],seed[2609],seed[644],seed[1602],seed[1230],seed[3919],seed[1044],seed[1264],seed[3181],seed[3982],seed[763],seed[443],seed[690],seed[1403],seed[1594],seed[1596],seed[2511],seed[1080],seed[759],seed[2260],seed[2120],seed[3246],seed[509],seed[2552],seed[3438],seed[3353],seed[899],seed[1812],seed[3770],seed[160],seed[3003],seed[3937],seed[336],seed[3200],seed[710],seed[822],seed[2165],seed[3754],seed[1549],seed[692],seed[3023],seed[3008],seed[528],seed[829],seed[3011],seed[2280],seed[394],seed[2322],seed[2123],seed[1540],seed[4044],seed[2300],seed[1752],seed[3822],seed[1418],seed[3032],seed[3990],seed[2801],seed[756],seed[2231],seed[133],seed[3009],seed[3431],seed[873],seed[3121],seed[1064],seed[1553],seed[1498],seed[3082],seed[454],seed[1480],seed[2833],seed[126],seed[2073],seed[2840],seed[516],seed[1245],seed[2004],seed[3598],seed[1010],seed[2628],seed[356],seed[874],seed[1682],seed[3680],seed[3541],seed[3306],seed[1558],seed[1804],seed[769],seed[1846],seed[3931],seed[3463],seed[2987],seed[3207],seed[1185],seed[2905],seed[1571],seed[196],seed[293],seed[309],seed[1788],seed[1445],seed[730],seed[705],seed[2638],seed[1244],seed[1197],seed[3382],seed[2561],seed[1489],seed[2002],seed[1255],seed[1588],seed[518],seed[1077],seed[1676],seed[1960],seed[2268],seed[2950],seed[435],seed[1022],seed[181],seed[4056],seed[172],seed[2025],seed[3604],seed[3649],seed[3543],seed[3544],seed[3869],seed[3445],seed[3000],seed[1680],seed[3467],seed[1743],seed[101],seed[1105],seed[1793],seed[3605],seed[918],seed[876],seed[307],seed[3566],seed[2528],seed[2171],seed[2645],seed[2388],seed[2730],seed[1236],seed[917],seed[3837],seed[642],seed[928],seed[4070],seed[3358],seed[1864],seed[3167],seed[2373],seed[436],seed[3153],seed[4064],seed[800],seed[3221],seed[3715],seed[746],seed[1569],seed[3917],seed[2124],seed[2575],seed[3711],seed[1668],seed[2410],seed[3086],seed[510],seed[3391],seed[2579],seed[2569],seed[3112],seed[3567],seed[1829],seed[2886],seed[3572],seed[408],seed[602],seed[494],seed[2078],seed[2360],seed[2199],seed[3944],seed[3069],seed[2145],seed[1740],seed[2258],seed[2877],seed[2968],seed[1707],seed[3089],seed[1645],seed[3460],seed[929],seed[3458],seed[213],seed[2254],seed[741],seed[2089],seed[270],seed[3847],seed[2847],seed[3122],seed[579],seed[69],seed[3994],seed[1981],seed[2719],seed[2342],seed[3385],seed[1275],seed[2924],seed[859],seed[3354],seed[3036],seed[2475],seed[3658],seed[3998],seed[2224],seed[4080],seed[473],seed[27],seed[1239],seed[2734],seed[1441],seed[2936],seed[2939],seed[0],seed[66],seed[2705],seed[2146],seed[3664],seed[666],seed[3712],seed[2928],seed[1938],seed[2027],seed[3969],seed[2181],seed[3141],seed[2602],seed[2327],seed[831],seed[30],seed[3224],seed[824],seed[983],seed[1739],seed[624],seed[3346],seed[87],seed[1593],seed[3550],seed[1231],seed[238],seed[227],seed[1665],seed[3893],seed[3643],seed[2088],seed[2084],seed[1550],seed[2862],seed[2346],seed[1714],seed[306],seed[206],seed[2899],seed[1263],seed[2396],seed[1590],seed[3242],seed[3925],seed[205],seed[3015],seed[1510],seed[2670],seed[3891],seed[2577],seed[3562],seed[95],seed[959],seed[839],seed[3345],seed[3046],seed[1268],seed[4003],seed[1127],seed[37],seed[244],seed[1867],seed[3007],seed[3648],seed[361],seed[1606],seed[3192],seed[290],seed[1206],seed[2625],seed[1822],seed[1880],seed[1116],seed[2681],seed[424],seed[1184],seed[3198],seed[3904],seed[486],seed[2518],seed[3965],seed[989],seed[177],seed[3555],seed[1333],seed[267],seed[531],seed[593],seed[1644],seed[2110],seed[312],seed[1546],seed[444],seed[1012],seed[2174],seed[1056],seed[2011],seed[1651],seed[1156],seed[2458],seed[2469],seed[2428],seed[695],seed[628],seed[536],seed[4085],seed[760],seed[1026],seed[1166],seed[366],seed[954],seed[1987],seed[3499],seed[1485],seed[1152],seed[3859],seed[1280],seed[320],seed[662],seed[1066],seed[2452],seed[4072],seed[1316],seed[977],seed[1218],seed[2026],seed[3582],seed[1209],seed[1154],seed[2588],seed[4008],seed[610],seed[1533],seed[682],seed[1327],seed[1384],seed[1774],seed[2777],seed[465],seed[3962],seed[2942],seed[1420],seed[3947],seed[527],seed[470],seed[2805],seed[2467],seed[2827],seed[1270],seed[41],seed[1934],seed[3208],seed[3481],seed[23],seed[114],seed[3935],seed[1458],seed[1642],seed[2385],seed[2715],seed[1059],seed[2824],seed[2739],seed[265],seed[1452],seed[1771],seed[1222],seed[1667],seed[3867],seed[341],seed[3180],seed[2901],seed[49],seed[2604],seed[3621],seed[1552],seed[2999],seed[1286],seed[3915],seed[2855],seed[3812],seed[251],seed[2434],seed[4083],seed[3482],seed[3154],seed[226],seed[2741],seed[2355],seed[3772],seed[3178],seed[3031],seed[4052],seed[2210],seed[1974],seed[2639],seed[1019],seed[936],seed[2230],seed[131],seed[1221],seed[2616],seed[3341],seed[1271],seed[2631],seed[2808],seed[1272],seed[310],seed[1990],seed[2857],seed[728],seed[3685],seed[1732],seed[693],seed[285],seed[890],seed[2724],seed[2269],seed[2876],seed[2606],seed[2894],seed[3357],seed[3166],seed[3209],seed[2851],seed[81],seed[604],seed[1611],seed[3150],seed[168],seed[333],seed[3229],seed[330],seed[167],seed[1702],seed[3101],seed[1337],seed[3104],seed[3188],seed[493],seed[1910],seed[452],seed[2885],seed[194],seed[1305],seed[2546],seed[4071],seed[2433],seed[1207],seed[3049],seed[1111],seed[3367],seed[3558],seed[3068],seed[2212],seed[153],seed[3570],seed[2585],seed[655],seed[346],seed[1917],seed[2223],seed[938],seed[3175],seed[76],seed[2315],seed[3421],seed[2214],seed[411],seed[1252],seed[354],seed[3173],seed[1748],seed[3284],seed[506],seed[3352],seed[2324],seed[2654],seed[2913],seed[3725],seed[1946],seed[337],seed[2105],seed[1138],seed[2108],seed[2063],seed[3073],seed[1005],seed[875],seed[2242],seed[3578],seed[3677],seed[236],seed[209],seed[340],seed[2232],seed[539],seed[900],seed[2972],seed[637],seed[1499],seed[2736],seed[317],seed[3155],seed[2170],seed[3136],seed[2157],seed[462],seed[2249],seed[382],seed[1970],seed[284],seed[269],seed[1781],seed[3797],seed[1210],seed[3940],seed[1400],seed[2997],seed[1963],seed[1520],seed[2557],seed[2096],seed[3312],seed[2062],seed[2679],seed[3678],seed[2465],seed[4074],seed[2257],seed[667],seed[15],seed[3355],seed[1158],seed[3608],seed[525],seed[3767],seed[3035],seed[2168],seed[2023],seed[2309],seed[201],seed[2295],seed[1455],seed[1741],seed[2226],seed[2633],seed[272],seed[1574],seed[659],seed[2772],seed[2329],seed[843],seed[3241],seed[1148],seed[53],seed[1758],seed[2485],seed[722],seed[798],seed[220],seed[453],seed[1],seed[1889],seed[944],seed[379],seed[1556],seed[198],seed[397],seed[2526],seed[908],seed[3879],seed[3957],seed[2237],seed[2816],seed[63],seed[86],seed[3138],seed[1841],seed[552],seed[1627],seed[3328],seed[3084],seed[2201],seed[975],seed[3875],seed[2412],seed[1968],seed[846],seed[3557],seed[3067],seed[2731],seed[3260],seed[127],seed[3507],seed[1634],seed[2795],seed[2982],seed[542],seed[3574],seed[2826],seed[1362],seed[119],seed[3790],seed[1411],seed[1899],seed[4067],seed[491],seed[3734],seed[2944],seed[1046],seed[1000],seed[3403],seed[1117],seed[1773],seed[274],seed[2172],seed[2319],seed[2314],seed[3014],seed[2690],seed[554],seed[3968],seed[2983],seed[3849],seed[994],seed[952],seed[1720],seed[3381],seed[384],seed[3936],seed[1211],seed[387],seed[35],seed[2325],seed[3816],seed[499],seed[3317],seed[3102],seed[568],seed[2044],seed[16],seed[249],seed[428],seed[3047],seed[3581],seed[1421],seed[2219],seed[3441],seed[386],seed[1199],seed[3446],seed[3363],seed[950],seed[943],seed[782],seed[605],seed[1028],seed[2523],seed[183],seed[2348],seed[3392],seed[2437],seed[2244],seed[3496],seed[3128],seed[3248],seed[3970],seed[322],seed[261],seed[180],seed[481],seed[74],seed[4001],seed[2185],seed[1967],seed[1195],seed[1192],seed[2184],seed[1332],seed[788],seed[3270],seed[2533],seed[3762],seed[3870],seed[1563],seed[1226],seed[1276],seed[3533],seed[4020],seed[749],seed[218],seed[4010],seed[3005],seed[2080],seed[862],seed[1399],seed[405],seed[1131],seed[1706],seed[3911],seed[2912],seed[417],seed[3475],seed[3537],seed[369],seed[1765],seed[3010],seed[3967],seed[3028],seed[2595],seed[1802],seed[1172],seed[3075],seed[4059],seed[371],seed[1145],seed[2299],seed[1745],seed[2411],seed[3587],seed[277],seed[2481],seed[479],seed[2574],seed[3662],seed[1531],seed[1323],seed[2720],seed[3286],seed[555],seed[3750],seed[2302],seed[3746],seed[3882],seed[3143],seed[2116],seed[821],seed[2748],seed[2821],seed[1352],seed[1512],seed[1129],seed[1496],seed[43],seed[2710],seed[1891],seed[2225],seed[2841],seed[4014],seed[1998],seed[3801],seed[264],seed[1360],seed[1173],seed[1081],seed[273],seed[1290],seed[3411],seed[399],seed[182],seed[651],seed[3930],seed[2043],seed[314],seed[999],seed[1777],seed[3806],seed[1959],seed[3855],seed[186],seed[3193],seed[857],seed[3251],seed[2275],seed[2854],seed[3182],seed[3996],seed[1047],seed[3839],seed[978],seed[2757],seed[968],seed[1054],seed[1536],seed[3730],seed[3227],seed[1449],seed[3512],seed[2618],seed[2147],seed[3300],seed[2284],seed[1826],seed[2454],seed[305],seed[2916],seed[378],seed[738],seed[2745],seed[2815],seed[3266],seed[2246],seed[1717],seed[1311],seed[3452],seed[1660],seed[3168],seed[3416],seed[2218],seed[3641],seed[3710],seed[3895],seed[1893],seed[3057],seed[1964],seed[2782],seed[3539],seed[1614],seed[94],seed[3199],seed[2006],seed[1196],seed[116],seed[4046],seed[3958],seed[2946],seed[3777],seed[4069],seed[3650],seed[1317],seed[3279],seed[3986],seed[2221],seed[629],seed[485],seed[2562],seed[3337],seed[2696],seed[2151],seed[1072],seed[2753],seed[2001],seed[1672],seed[401],seed[221],seed[764],seed[3447],seed[3657],seed[2473],seed[2769],seed[5],seed[2883],seed[2892],seed[1730],seed[3485],seed[2358],seed[735],seed[3589],seed[1457],seed[3955],seed[2176],seed[3542],seed[197],seed[1204],seed[1969],seed[1374],seed[2292],seed[3984],seed[627],seed[577],seed[3766],seed[316],seed[3681],seed[2903],seed[1477],seed[1393],seed[2138],seed[3090],seed[4051],seed[2182],seed[2103],seed[2694],seed[1709],seed[2444],seed[1671],seed[2127],seed[3885],seed[3486],seed[2713],seed[2251],seed[1798],seed[3360],seed[988],seed[159],seed[926],seed[3034],seed[849],seed[2861],seed[4049],seed[2553],seed[476],seed[2156],seed[573],seed[145],seed[304],seed[3051],seed[956],seed[704],seed[174],seed[1159],seed[1902],seed[3577],seed[1699],seed[920],seed[911],seed[1067],seed[1168],seed[3756],seed[1112],seed[255],seed[622],seed[2441],seed[1681],seed[1342],seed[3894],seed[3856],seed[105],seed[1189],seed[3302],seed[2943],seed[3946],seed[2404],seed[2989],seed[565],seed[699],seed[923],seed[263],seed[1643],seed[3272],seed[2197],seed[1139],seed[2525],seed[3097],seed[1492],seed[3659],seed[1467],seed[670],seed[1823],seed[634],seed[1101],seed[191],seed[1381],seed[3289],seed[2427],seed[3281],seed[3440],seed[3303],seed[1750],seed[2440],seed[2693],seed[1238],seed[3370],seed[2093],seed[884],seed[773],seed[784],seed[3732],seed[78],seed[3778],seed[1202],seed[1971],seed[3961],seed[179],seed[3022],seed[297],seed[2934],seed[2742],seed[1795],seed[684],seed[2935],seed[2457],seed[2798],seed[2049],seed[903],seed[18],seed[3860],seed[1504],seed[1723],seed[2991],seed[1309],seed[2099],seed[3615],seed[3943],seed[1205],seed[3886],seed[3085],seed[2399],seed[2464],seed[2126],seed[797],seed[1090],seed[3245],seed[2121],seed[146],seed[3887],seed[976],seed[115],seed[861],seed[2035],seed[955],seed[1338],seed[614],seed[3497],seed[2367],seed[1843],seed[1888],seed[1876],seed[1575],seed[3335],seed[1383],seed[1208],seed[1216],seed[3350],seed[1108],seed[1503],seed[3724],seed[3872],seed[294],seed[836],seed[706],seed[2010],seed[1160],seed[3479],seed[2304],seed[790],seed[1017],seed[440],seed[4057],seed[2548],seed[474],seed[582],seed[2328],seed[2783],seed[3186],seed[2175],seed[1014],seed[2293],seed[1701],seed[887],seed[3989],seed[2253],seed[2867],seed[1137],seed[2990],seed[3118],seed[3261],seed[1578],seed[2613],seed[1475],seed[649],seed[2590],seed[656],seed[827],seed[1435],seed[1490],seed[1919],seed[353],seed[3201],seed[1863],seed[2177],seed[2965],seed[3393],seed[3742],seed[775],seed[2429],seed[1735],seed[1976],seed[2270],seed[1120],seed[325],seed[592],seed[3365],seed[916],seed[2592],seed[647],seed[2298],seed[3857],seed[2586],seed[894],seed[1494],seed[47],seed[2104],seed[2708],seed[2929],seed[3383],seed[162],seed[1165],seed[2289],seed[3030],seed[433],seed[4025],seed[323],seed[1178],seed[3442],seed[1821],seed[276],seed[4058],seed[1769],seed[740],seed[2305],seed[4030],seed[3660],seed[3796],seed[1083],seed[2608],seed[2852],seed[2770],seed[743],seed[3607],seed[1417],seed[36],seed[202],seed[3202],seed[2220],seed[3269],seed[1087],seed[268],seed[707],seed[1171],seed[2597],seed[92],seed[2800],seed[1235],seed[638],seed[1355],seed[472],seed[772],seed[501],seed[224],seed[1977],seed[3980],seed[1591],seed[946],seed[3709],seed[2313],seed[3928],seed[2276],seed[3080],seed[4043],seed[1647],seed[1240],seed[2067],seed[62],seed[1772],seed[3686],seed[2066],seed[3890],seed[2976],seed[1625],seed[144],seed[2317],seed[2306],seed[3902],seed[3617],seed[1203],seed[3819],seed[3361],seed[135],seed[67],seed[2986],seed[583],seed[79],seed[2310],seed[3956],seed[3752],seed[3760],seed[3025],seed[3287],seed[2308],seed[818],seed[2507],seed[2765],seed[2759],seed[2729],seed[2352],seed[2274],seed[1088],seed[3165],seed[1537],seed[2402],seed[2476],seed[2530],seed[3521],seed[381],seed[2278],seed[3],seed[3152],seed[3763],seed[3206],seed[2637],seed[3222],seed[2674],seed[538],seed[1057],seed[3735],seed[3805],seed[260],seed[2071],seed[3765],seed[567],seed[3802],seed[3768],seed[2107],seed[1678],seed[3726],seed[3111],seed[3784],seed[10],seed[2911],seed[2227],seed[2233],seed[2871],seed[231],seed[1903],seed[3119],seed[1130],seed[2921],seed[3472],seed[2144],seed[3861],seed[3618],seed[1652],seed[3487],seed[2164],seed[2747],seed[1937],seed[2763],seed[2682],seed[3842],seed[598],seed[3716],seed[2996],seed[2020],seed[2417],seed[1636],seed[1307],seed[3653],seed[2688],seed[3776],seed[1605],seed[3788],seed[111],seed[3545],seed[674],seed[3336],seed[3547],seed[3863],seed[1147],seed[451],seed[1291],seed[1434],seed[3780],seed[985],seed[2413],seed[505],seed[522],seed[364],seed[1308],seed[3164],seed[3978],seed[4036],seed[2393],seed[3058],seed[2834],seed[632],seed[3810],seed[3525],seed[1713],seed[2593],seed[913],seed[2450],seed[3783],seed[2646],seed[2802],seed[1901],seed[2610],seed[2259],seed[2432],seed[2790],seed[3723],seed[166],seed[1297],seed[2909],seed[2754],seed[3546],seed[3619],seed[1016],seed[912],seed[1710],seed[981],seed[3439],seed[1414],seed[2543],seed[1190],seed[925],seed[816],seed[243],seed[2055],seed[825],seed[4031],seed[1658],seed[123],seed[3912],seed[686],seed[45],seed[2522],seed[82],seed[219],seed[2860],seed[558],seed[2390],seed[940],seed[217],seed[332],seed[1554],seed[3390],seed[1508],seed[1613],seed[3927],seed[3278],seed[138],seed[2069],seed[1965],seed[3285],seed[963],seed[4005],seed[3434],seed[2849],seed[3817],seed[2621],seed[90],seed[3437],seed[2125],seed[2262],seed[377],seed[2200],seed[3296],seed[2050],seed[4000],seed[132],seed[3596],seed[1657],seed[4093],seed[3744],seed[2307],seed[2953],seed[2162],seed[3637],seed[2247],seed[3157],seed[1814],seed[24],seed[708],seed[2704],seed[1181],seed[2836],seed[1993],seed[3921],seed[59],seed[4055],seed[1033],seed[1128],seed[3065],seed[2799],seed[2158],seed[3459],seed[2409],seed[1320],seed[1945],seed[2650],seed[3652],seed[3638],seed[4012],seed[1753],seed[2607],seed[1683],seed[612],seed[3140],seed[543],seed[3484],seed[1514],seed[524],seed[2531],seed[2668],seed[1861],seed[1187],seed[609],seed[1346],seed[1126],seed[2947],seed[1053],seed[2179],seed[3673],seed[3597],seed[1906],seed[712],seed[1687],seed[3061],seed[530],seed[19],seed[2766],seed[3282],seed[2920],seed[3430],seed[2949],seed[1348],seed[844],seed[1201],seed[838],seed[2029],seed[2466],seed[1925],seed[3888],seed[3339],seed[2436],seed[455],seed[553],seed[1365],seed[1640],seed[1896],seed[1905],seed[1871],seed[3883],seed[2534],seed[2418],seed[3062],seed[1132],seed[3257],seed[1862],seed[3899],seed[3076],seed[2395],seed[52],seed[3462],seed[1102],seed[3158],seed[3571],seed[3683],seed[1283],seed[1689],seed[3183],seed[1227],seed[2647],seed[3833],seed[288],seed[747],seed[2122],seed[2829],seed[2738],seed[1432],seed[3591],seed[2699],seed[3056],seed[2890],seed[3593],seed[2510],seed[2297],seed[1106],seed[2282],seed[2456],seed[477],seed[3297],seed[2728],seed[345],seed[2271],seed[3029],seed[3457],seed[2767],seed[1061],seed[1140],seed[107],seed[3268],seed[3351],seed[289],seed[100],seed[930],seed[678],seed[2888],seed[88],seed[1279],seed[1464],seed[2709],seed[1186],seed[1161],seed[2167],seed[1143],seed[3914],seed[2971],seed[3654],seed[2128],seed[2975],seed[1935],seed[2505],seed[3785],seed[1078],seed[2028],seed[1724],seed[91],seed[3469],seed[1560],seed[3079],seed[2814],seed[2707],seed[315],seed[414],seed[3612],seed[3506],seed[860],seed[1956],seed[3749],seed[1595],seed[1095],seed[1736],seed[786],seed[338],seed[56],seed[2420],seed[902],seed[504],seed[129],seed[3362],seed[1242],seed[3397],seed[1448],seed[2111],seed[3731],seed[2733],seed[4090],seed[2149],seed[3556],seed[3689],seed[1799],seed[2740],seed[1409],seed[2558],seed[1879],seed[1887],seed[2286],seed[3532],seed[2141],seed[1287],seed[3616],seed[1587],seed[939],seed[3705],seed[3694],seed[702],seed[2915],seed[42],seed[1326],seed[3908],seed[1356],seed[223],seed[868],seed[2686],seed[3418],seed[3324],seed[4065],seed[204],seed[2132],seed[2488],seed[2662],seed[2007],seed[2692],seed[1113],seed[1426],seed[3600],seed[3864],seed[12],seed[2596],seed[70],seed[2046],seed[3332],seed[2135],seed[636],seed[980],seed[2098],seed[3918],seed[619],seed[2204],seed[1149],seed[390],seed[1986],seed[3410],seed[1405],seed[2567],seed[1616],seed[2508],seed[3117],seed[3661],seed[1727],seed[1661],seed[3059],seed[3255],seed[533],seed[2323],seed[502],seed[2446],seed[3129],seed[842],seed[1872],seed[2169],seed[1921],seed[1382],seed[2619],seed[2287],seed[1366],seed[2906],seed[3413],seed[576],seed[3929],seed[1979],seed[1465],seed[3502],seed[1809],seed[3432],seed[3323],seed[2605],seed[2573],seed[357],seed[630],seed[3798],seed[3540],seed[427],seed[2572],seed[1371],seed[669],seed[2524],seed[3233],seed[1251],seed[2261],seed[407],seed[3877],seed[4013],seed[723],seed[2166],seed[854],seed[635],seed[3223],seed[3687],seed[2474],seed[256],seed[1237],seed[1629],seed[1631],seed[834],seed[3012],seed[1786],seed[1819],seed[2335],seed[1856],seed[3315],seed[134],seed[1328],seed[2559],seed[3625],seed[4039],seed[886],seed[713],seed[1731],seed[2615],seed[1599],seed[1091],seed[318],seed[3960],seed[410],seed[2114],seed[1122],seed[2130],seed[3874],seed[1573],seed[863],seed[3124],seed[2571],seed[2239],seed[450],seed[785],seed[4],seed[3713],seed[3519],seed[965],seed[3628],seed[239],seed[2865],seed[1150],seed[3633],seed[673],seed[2891],seed[2431],seed[2015],seed[120],seed[2374],seed[1991],seed[2497],seed[663],seed[2058],seed[1547],seed[334],seed[3103],seed[233],seed[2653],seed[2490],seed[828],seed[648],seed[896],seed[3349],seed[1583],seed[789],seed[3375],seed[3120],seed[3342],seed[534],seed[3741],seed[3682],seed[383],seed[2514],seed[3037],seed[645],seed[3108],seed[3247],seed[2962],seed[1598],seed[2599],seed[3088],seed[3169],seed[1927],seed[3624],seed[1722],seed[208],seed[1422],seed[1153],seed[3027],seed[2148],seed[1728],seed[1637],seed[3516],seed[1110],seed[1559],seed[3923],seed[2846],seed[588],seed[4092],seed[570],seed[2521],seed[3275],seed[2520],seed[199],seed[2551],seed[2192],seed[1146],seed[556],seed[1674],seed[744],seed[2294],seed[3074],seed[1104],seed[2835],seed[1258],seed[388],seed[979],seed[545],seed[1663],seed[2252],seed[2318],seed[719],seed[2874],seed[4073],seed[2687],seed[3853],seed[3004],seed[3319],seed[2830],seed[280],seed[1200],seed[2651],seed[1176],seed[38],seed[185],seed[3376],seed[3477],seed[1483],seed[2248],seed[2109],seed[1865],seed[858],seed[4045],seed[3811],seed[3053],seed[1357],seed[660],seed[3288],seed[2459],seed[3603],seed[2034],seed[1164],seed[2760],seed[2701],seed[1797],seed[914],seed[3252],seed[4076],seed[2052],seed[235],seed[2316],seed[3972],seed[1949],seed[3913],seed[2054],seed[1783],seed[599],seed[3399],seed[3114],seed[99],seed[1314],seed[847],seed[2914],seed[3561],seed[3708],seed[1516],seed[490],seed[2718],seed[17],seed[595],seed[701],seed[26],seed[1923],seed[2414],seed[1368],seed[2353],seed[3953],seed[1827],seed[2272],seed[3283],seed[3954],seed[757],seed[953],seed[561],seed[178],seed[1733],seed[3535],seed[2356],seed[3292],seed[61],seed[574],seed[1519],seed[2372],seed[3271],seed[590],seed[1794],seed[2664],seed[1756],seed[3718],seed[3344],seed[1911],seed[1789],seed[1751],seed[1719],seed[3728],seed[3588],seed[1900],seed[2797],seed[724],seed[1438],seed[4075],seed[475],seed[3425],seed[1300],seed[681],seed[813],seed[3256],seed[2207],seed[1757],seed[2758],seed[3017],seed[3389],seed[3523],seed[1339],seed[3396],seed[520],seed[136],seed[1768],seed[3348],seed[3733],seed[3013],seed[3384],seed[1858],seed[1424],seed[2764],seed[2375],seed[2925],seed[2931],seed[1655],seed[1466],seed[3629],seed[2076],seed[1749],seed[148],seed[3951],seed[1032],seed[426],seed[2471],seed[34],seed[2667],seed[3039],seed[2630],seed[537],seed[2101],seed[1386],seed[2256],seed[594],seed[4053],seed[3636],seed[375],seed[1479],seed[1632],seed[1505],seed[3826],seed[1961],seed[1646],seed[2863],seed[1299],seed[229],seed[3455],seed[855],seed[2509],seed[780],seed[616],seed[1779],seed[3721],seed[2695],seed[1040],seed[1407],seed[3920],seed[626],seed[319],seed[871],seed[164],seed[2008],seed[3042],seed[1058],seed[3020],seed[2979],seed[3041],seed[3906],seed[1350],seed[984],seed[2542],seed[3809],seed[951],seed[2243],seed[889],seed[1079],seed[734],seed[3670],seed[2478],seed[3676],seed[3568],seed[3184],seed[3595],seed[3083],seed[434],seed[275],seed[1851],seed[4009],seed[819],seed[736],seed[3758],seed[3774],seed[1952],seed[1897],seed[2153],seed[1633],seed[2545],seed[3761],seed[3449],seed[907],seed[1524],seed[2194],seed[2967],seed[549],seed[2649],seed[1343],seed[2344],seed[1228],seed[2685],seed[1972],seed[1545],seed[2266],seed[3294],seed[2658],seed[809],seed[2094],seed[2363],seed[1796],seed[3702],seed[2455],seed[1468],seed[3189],seed[1572],seed[2584],seed[2462],seed[142],seed[812],seed[1517],seed[2812],seed[814],seed[1840],seed[1018],seed[2461],seed[3696],seed[3706],seed[1580],seed[503],seed[1764],seed[802],seed[1626],seed[1315],seed[2143],seed[3379],seed[2952],seed[2406],seed[2671],seed[3318],seed[3747],seed[2235],seed[3828],seed[3264],seed[1369],seed[3854],seed[1493],seed[3720],seed[3808],seed[1020],seed[3087],seed[1260],seed[3021],seed[3795],seed[1319],seed[328],seed[2351],seed[877],seed[1568],seed[3018],seed[1335],seed[1985],seed[1557],seed[2722],seed[193],seed[498],seed[3427],seed[2228],seed[600],seed[2850],seed[3064],seed[1778],seed[207],seed[363],seed[449],seed[3215],seed[4048],seed[1246],seed[1914],seed[4027],seed[3896],seed[4023],seed[413],seed[2036],seed[562],seed[1313],seed[2743],seed[2097],seed[1695],seed[141],seed[3668],seed[966],seed[33],seed[1141],seed[2350],seed[1834],seed[3259],seed[737],seed[2828],seed[547],seed[1274],seed[2768],seed[2453],seed[3214],seed[2477],seed[883],seed[3719],seed[2908],seed[1780],seed[1673],seed[29],seed[2540],seed[3693],seed[3498],seed[1004],seed[3737],seed[2755],seed[2676],seed[1446],seed[484],seed[1922],seed[3038],seed[339],seed[792],seed[2697],seed[4091],seed[2794],seed[3408],seed[3395],seed[535],seed[3775],seed[3078],seed[1878],seed[3356],seed[1530],seed[2236],seed[3309],seed[526],seed[841],seed[2725],seed[650],seed[3197],seed[3821],seed[2472],seed[2095],seed[687],seed[1670],seed[2726],seed[658],seed[948],seed[575],seed[3916],seed[2493],seed[2938],seed[2030],seed[2875],seed[4029],seed[3422],seed[3889],seed[3273],seed[1742],seed[3131],seed[222],seed[2019],seed[3474],seed[3634],seed[2386],seed[1125],seed[3651],seed[3156],seed[927],seed[606],seed[2555],seed[941],seed[2869],seed[3398],seed[1828],seed[1607],seed[2864],seed[1296],seed[905],seed[1940],seed[2154],seed[3196],seed[2354],seed[3979],seed[303],seed[3443],seed[1292],seed[1423],seed[4034],seed[3580],seed[3552],seed[2910],seed[2403],seed[4032],seed[1784],seed[1071],seed[327],seed[3132],seed[3663],seed[2012],seed[1413],seed[3448],seed[1182],seed[3941],seed[3191],seed[3602],seed[3254],seed[329],seed[2378],seed[2070],seed[1213],seed[3126],seed[1712],seed[3170],seed[3220],seed[717],seed[910],seed[2504],seed[1249],seed[3490],seed[691],seed[3262],seed[3656],seed[1523],seed[237],seed[1609],seed[837],seed[1581],seed[1838],seed[1043],seed[2749],seed[1877],seed[3782],seed[1837],seed[1930],seed[1694],seed[3428],seed[2330],seed[3583],seed[1388],seed[487],seed[1170],seed[2626],seed[869],seed[2326],seed[2032],seed[1848],seed[2479],seed[171],seed[2113],seed[1391],seed[348],seed[2882],seed[1617],seed[3697],seed[175],seed[1770],seed[3831],seed[897],seed[2907],seed[28],seed[1135],seed[3423],seed[102],seed[731],seed[2784],seed[2380],seed[2970],seed[2904],seed[1015],seed[3692],seed[1918],seed[2617],seed[2206],seed[402],seed[2632],seed[1100],seed[803],seed[165],seed[1886],seed[2727],seed[853],seed[3293],seed[685],seed[2347],seed[3844],seed[2215],seed[1076],seed[124],seed[1118],seed[720],seed[415],seed[508],seed[1615],seed[3301],seed[1261],seed[4007],seed[3959],seed[3703],seed[2640],seed[2536],seed[2622],seed[895],seed[1544],seed[40],seed[1232],seed[1373],seed[2312],seed[98],seed[935],seed[254],seed[1853],seed[1939],seed[2778],seed[3135],seed[3530],seed[832],seed[721],seed[3380],seed[2336],seed[431],seed[3372],seed[77],seed[2415],seed[1608],seed[3401],seed[3868],seed[480],seed[1041],seed[1295],seed[3331],seed[152],seed[711],seed[1639],seed[72],seed[960],seed[2387],seed[3509],seed[845],seed[3992],seed[2995],seed[970],seed[3926],seed[3225],seed[1395],seed[3415],seed[2423],seed[4033],seed[2937],seed[901],seed[1589],seed[3195],seed[1324],seed[3977],seed[2240],seed[3579],seed[1577],seed[1996],seed[3609],seed[1570],seed[1535],seed[2872],seed[3901],seed[810],seed[4060],seed[75],seed[932],seed[3329],seed[625],seed[856],seed[2222],seed[2343],seed[2059],seed[3759],seed[1430],seed[2974],seed[460],seed[2405],seed[2661],seed[4002],seed[1664],seed[2408],seed[416],seed[1055],seed[1436],seed[389],seed[3304],seed[3123],seed[2998],seed[1501],seed[3263],seed[4087],seed[3938],seed[2443],seed[2340],seed[1298],seed[1542],seed[794],seed[380],seed[1488],seed[1656],seed[548],seed[1451],seed[1973],seed[2893],seed[640],seed[3134],seed[3932],seed[3613],seed[2416],seed[3518],seed[1217],seed[3127],seed[343],seed[540],seed[2837],seed[2048],seed[257],seed[3404],seed[302],seed[65],seed[804],seed[1119],seed[2484],seed[3818],seed[2988],seed[2022],seed[1481],seed[489],seed[3374],seed[2897],seed[1364],seed[2021],seed[2535],seed[992],seed[1269],seed[2956],seed[993],seed[1460],seed[1994],seed[3646],seed[3834],seed[1321],seed[441],seed[1404],seed[2039],seed[791],seed[103],seed[3113],seed[3995],seed[362],seed[2072],seed[3631],seed[311],seed[3517],seed[2460],seed[3274],seed[1932],seed[2657],seed[891],seed[446],seed[1392],seed[3205],seed[3966],seed[1500],seed[3569],seed[3876],seed[2499],seed[1708],seed[1836],seed[1690],seed[2933],seed[32],seed[2680],seed[866],seed[1686],seed[2684],seed[513],seed[2161],seed[3866],seed[2614],seed[1134],seed[3063],seed[517],seed[921],seed[3298],seed[1995],seed[2005],seed[1476],seed[3325],seed[2842],seed[3804],seed[3414],seed[3204],seed[97],seed[1486],seed[922],seed[3240],seed[1233],seed[117],seed[1803],seed[807],seed[3492],seed[3310],seed[709],seed[2320],seed[1484],seed[2873],seed[1805],seed[2321],seed[2364],seed[1954],seed[1926],seed[1532],seed[4095],seed[2537],seed[3016],seed[727],seed[1459],seed[1241],seed[2868],seed[4068],seed[2856],seed[1285],seed[430],seed[1635],seed[2018],seed[621],seed[2969],seed[2234],seed[661],seed[2376],seed[1820],seed[945],seed[3865],seed[2425],seed[1303],seed[1624],seed[2331],seed[3420],seed[2024],seed[2000],seed[739],seed[1791],seed[3322],seed[1641],seed[283],seed[3534],seed[3549],seed[1738],seed[1390],seed[1062],seed[1450],seed[1539],seed[187],seed[2337],seed[1763],seed[1385],seed[406],seed[958],seed[2663],seed[688],seed[551],seed[2160],seed[2397],seed[589],seed[372],seed[1021],seed[1978],seed[689],seed[39],seed[2918],seed[55],seed[1497],seed[3513],seed[2612],seed[11],seed[2641],seed[677],seed[1329],seed[3983],seed[3666],seed[1097],seed[21],seed[3942],seed[1225],seed[301],seed[1243],seed[3105],seed[2419],seed[1431],seed[2196],seed[3444],seed[1666],seed[1868],seed[2051],seed[1133],seed[463],seed[3489],seed[808],seed[1928],seed[4088],seed[1529],seed[3308],seed[292],seed[2756],seed[425],seed[2655],seed[698],seed[1439],seed[633],seed[3655],seed[1412],seed[1920],seed[2487],seed[149],seed[2213],seed[93],seed[1885],seed[211],seed[2085],seed[3559],seed[3066],seed[1157],seed[2624],seed[266],seed[2566],seed[1792],seed[1755],seed[982],seed[4089],seed[7],seed[2642],seed[1693],seed[1725],seed[2838],seed[1001],seed[1654],seed[2065],seed[3473],seed[3213],seed[1705],seed[2702],seed[1194],seed[783],seed[1094],seed[2277],seed[1951],seed[157],seed[885],seed[1600],seed[3216],seed[3321],seed[1844],seed[3077],seed[2332],seed[3647],seed[2057],seed[1565],seed[833],seed[3386],seed[3779],seed[3433],seed[3903],seed[2635],seed[1815],seed[2594],seed[2656],seed[665],seed[541],seed[3727],seed[3584],seed[3755],seed[3508],seed[4079],seed[3878],seed[3981],seed[615],seed[664],seed[766],seed[1254],seed[3642],seed[271],seed[2470],seed[3226],seed[3159],seed[1869],seed[1188],seed[779],seed[733],seed[2383],seed[942],seed[2482],seed[3851],seed[3799],seed[801],seed[3910],seed[2163],seed[3846],seed[618],seed[467],seed[3424],seed[3892],seed[2698],seed[1831],seed[512],seed[2880],seed[3050],seed[1267],seed[585],seed[3820],seed[3234],seed[3852],seed[3740],seed[3585],seed[872],seed[1331],seed[203],seed[557],seed[6],seed[1966],seed[3950],seed[2993],seed[3160],seed[2042],seed[1376],seed[31],seed[110],seed[1253],seed[3684],seed[195],seed[1069],seed[820],seed[287],seed[795],seed[1622],seed[13],seed[421],seed[3369],seed[3291],seed[2279],seed[671],seed[3897],seed[971],seed[3095],seed[987],seed[2819],seed[4037],seed[3092],seed[1312],seed[1334],seed[2463],seed[3040],seed[1944],seed[3531],seed[1669],seed[3503],seed[1592],seed[2014],seed[3594],seed[458],seed[3526],seed[776],seed[1304],seed[1857],seed[365],seed[2371],seed[2538],seed[1787],seed[478],seed[3945],seed[1515],seed[358],seed[796],seed[2980],seed[2775],seed[1782],seed[2576],seed[1219],seed[3840],seed[459],seed[3949],seed[3099],seed[3149],seed[3347],seed[1419],seed[2291],seed[2807],seed[2583],seed[3807],seed[2737],seed[4086],seed[683],seed[563],seed[1220],seed[3622],seed[2091],seed[2361],seed[1845],seed[2515],seed[4042],seed[2940],seed[176],seed[514],seed[2031],seed[2627],seed[1586],seed[2564],seed[4015],seed[3773],seed[623],seed[1566],seed[1543],seed[423],seed[497],seed[3674],seed[2117],seed[2193],seed[1754],seed[2879],seed[2480],seed[560],seed[1638],seed[1082],seed[3501],seed[3054],seed[300],seed[1847],seed[3144],seed[2691],seed[3212],seed[2550],seed[2195],seed[1527],seed[781],seed[3453],seed[4016],seed[121],seed[2392],seed[793],seed[753],seed[1433],seed[2496],seed[1175],seed[2285],seed[591],seed[1711],seed[3743],seed[212],seed[1103],seed[360],seed[3825],seed[4061],seed[2498],seed[1953],seed[750],seed[2957],seed[2889],seed[1256],seed[3769],seed[3880],seed[3848],seed[216],seed[1471],seed[1620],seed[3898],seed[2845],seed[2881],seed[3190],seed[1347],seed[1401],seed[1833],seed[3841],seed[2774],seed[4019],seed[1415],seed[694],seed[2506],seed[1049],seed[3174],seed[2930],seed[1759],seed[2366],seed[3794],seed[1470],seed[214],seed[404],seed[777],seed[3873],seed[1367],seed[3973],seed[3468],seed[242],seed[3265],seed[1507],seed[654],seed[3177],seed[409],seed[1025],seed[22],seed[986],seed[607],seed[1406],seed[3176],seed[2438],seed[2365],seed[104],seed[2791],seed[2750],seed[2083],seed[48],seed[225],seed[1692],seed[787],seed[2955],seed[1281],seed[3280],seed[3757],seed[3081],seed[3627],seed[3738],seed[3239],seed[1904],seed[2926],seed[3210],seed[3388],seed[3172],seed[1700],seed[2703],seed[2037],seed[1474],seed[1734],seed[1289],seed[1518],seed[2381],seed[1999],seed[1988],seed[1950],seed[2611],seed[597],seed[3464],seed[3748],seed[96],seed[3217],seed[1068],seed[1003],seed[1597],seed[973],seed[3522],seed[246],seed[878],seed[278],seed[904],seed[2789],seed[2665],seed[3002],seed[3753],seed[370],seed[2136],seed[393],seed[2424],seed[1525],seed[2556],seed[438],seed[1379],seed[113],seed[1548],seed[934],seed[3704],seed[2502],seed[1648],seed[1808],seed[1051],seed[2301],seed[758],seed[2217],seed[3793],seed[1807],seed[3070],seed[937],seed[2721],seed[2013],seed[2866],seed[725],seed[3491],seed[3644],seed[1506],seed[1013],seed[4035],seed[3871],seed[1612],seed[2963],seed[240],seed[20],seed[1601],seed[3564],seed[3402],seed[933],seed[3900],seed[1567],seed[1098],seed[1721],seed[2648],seed[385],seed[2486],seed[3480],seed[774],seed[3739],seed[2339],seed[3515],seed[1322],seed[3218],seed[2853],seed[2932],seed[2255],seed[2673],seed[752],seed[188],seed[1375],seed[58],seed[1060],seed[3368],seed[73],seed[147],seed[3707],seed[639],seed[1582],seed[326],seed[4081],seed[230],seed[2981],seed[2512],seed[445],seed[471],seed[4066],seed[2483],seed[2820],seed[3639],seed[299],seed[3466],seed[3091],seed[2563],seed[2539],seed[1163],seed[715],seed[308],seed[184],seed[2554],seed[569],seed[2400],seed[2825],seed[1907],seed[1746],seed[2549],seed[64],seed[51],seed[1027],seed[2785],seed[3745],seed[566],seed[2439],seed[190],seed[1183],seed[2643],seed[4028],seed[601],seed[466],seed[995],seed[3791],seed[2964],seed[2090],seed[3700],seed[2303],seed[2449],seed[2818],seed[2033],seed[68],seed[2788],seed[2810],seed[2341],seed[2263],seed[1358],seed[2142],seed[2283],seed[2370],seed[1007],seed[1943],seed[464],seed[3451],seed[716],seed[3044],seed[1982],seed[352],seed[2190],seed[2919],seed[2858],seed[2045],seed[295],seed[2202],seed[2811],seed[3614],seed[2448],seed[3813],seed[2009],seed[3026],seed[2334],seed[1980],seed[432],seed[1957],seed[2848],seed[703],seed[3277],seed[3417],seed[2809],seed[3109],seed[335],seed[578],seed[2839],seed[1234],seed[1958],seed[3688],seed[1619],seed[1491],seed[3714],seed[652],seed[2081],seed[2659],seed[1302],seed[2532],seed[1114],seed[3884],seed[3907],seed[3536],seed[3258],seed[2369],seed[1551],seed[2744],seed[961],seed[1775],seed[1093],seed[1810],seed[2112],seed[3244],seed[2500],seed[439],seed[653],seed[962],seed[4094],seed[1282],seed[1398],seed[3554],seed[3771],seed[1801],seed[1073],seed[1850],seed[2152],seed[3905],seed[2859],seed[852],seed[2951],seed[3789],seed[1852],seed[1354],seed[1402],seed[3985],seed[2394],seed[1817],seed[2115],seed[1790],seed[3729],seed[2106],seed[2422],seed[1036],seed[150],seed[2973],seed[2273],seed[2064],seed[521],seed[2706],seed[919],seed[641],seed[2016],seed[3881],seed[2541],seed[2519],seed[192],seed[3699],seed[1229],seed[1045],seed[2844],seed[2079],seed[130],seed[546],seed[44],seed[1691],seed[2945],seed[2100],seed[3148],seed[1151],seed[3326],seed[3232],seed[4054],seed[1830],seed[2779],seed[2389],seed[2773],seed[3161],seed[830],seed[2155],seed[2634],seed[696],seed[2966],seed[1121],seed[321],seed[515],seed[550],seed[3314],seed[3320],seed[2178],seed[1248],seed[879],seed[1169],seed[2384],seed[1716],seed[732],seed[3832],seed[1955],seed[1942],seed[949],seed[3922],seed[1881],seed[1854],seed[3429],seed[2205],seed[2445],seed[668],seed[584],seed[1340],seed[1469],seed[646],seed[2],seed[1265],seed[586],seed[3024],seed[2345],seed[2513],seed[8],seed[437],seed[2762],seed[882],seed[1380],seed[108],seed[2265],seed[3999],seed[1806],seed[2752],seed[1191],seed[1009],seed[1344],seed[751],seed[3470],seed[679],seed[2435],seed[398],seed[3231],seed[3338],seed[2985],seed[1992],seed[867],seed[2652],seed[1447],seed[3601],seed[400],seed[2771],seed[2296],seed[2817],seed[3611],seed[2229],seed[3514],seed[3052],seed[1038],seed[210],seed[1325],seed[3988],seed[2060],seed[3667],seed[2560],seed[1704],seed[3575],seed[457],seed[1223],seed[2250],seed[109],seed[3691],seed[1534],seed[2264],seed[523],seed[1099],seed[140],seed[2077],seed[54],seed[2187],seed[3290],seed[697],seed[1762],seed[3645],seed[392],seed[865],seed[2994],seed[1875],seed[241],seed[1330],seed[291],seed[3203],seed[3800],seed[906],seed[3630],seed[2047],seed[14],seed[888],seed[3909],seed[3327],seed[544],seed[3476],seed[3316],seed[1618],seed[1747],seed[2150],seed[158],seed[1277],seed[2732],seed[3071],seed[1372],seed[2672],seed[3493],seed[1662],seed[2430],seed[532],seed[247],seed[1924],seed[3299],seed[2407],seed[1389],seed[2186],seed[2377],seed[1603],seed[3100],seed[3243],seed[3751],seed[1039],seed[4022],seed[3520],seed[2338],seed[1425],seed[331],seed[745],seed[2129],seed[1528],seed[998],seed[3836],seed[3048],seed[447],seed[3426],seed[2442],seed[3971],seed[1306],seed[1034],seed[1895],seed[997],seed[1361],seed[915],seed[2191],seed[3238],seed[422],seed[374],seed[2600],seed[1074],seed[811],seed[2978],seed[373],seed[3764],seed[3933],seed[2644],seed[3675],seed[3610],seed[3671],seed[488],seed[1050],seed[342],seed[3378],seed[2238],seed[2580],seed[2677],seed[817],seed[3359],seed[3006],seed[3093],seed[1744],seed[350],seed[765],seed[3505],seed[2501],seed[1933],seed[3219],seed[611],seed[57],seed[3060],seed[2211],seed[1948],seed[1084],seed[3276],seed[420],seed[469],seed[893],seed[3620],seed[1684],seed[1541],seed[169],seed[1698],seed[1818],seed[1262],seed[2780],seed[344],seed[2902],seed[2581],seed[2620],seed[84],seed[3511],seed[1224],seed[2492],seed[3529],seed[1538],seed[3843],seed[3249],seed[3435],seed[840],seed[2717],seed[3151],seed[2139],seed[351],seed[3236],seed[1884],seed[83],seed[1679],seed[2751],seed[3098],seed[3137],seed[2675],seed[2578],seed[2603],seed[4041],seed[2714],seed[1162],seed[2636],seed[1284],seed[395],seed[419],seed[1177],seed[3106],seed[2958],seed[2568],seed[1011],seed[1048],seed[3551],seed[2203],seed[2491],seed[2922],seed[3538],seed[1136],seed[1070],seed[1677],seed[1456],seed[2041],seed[1630],seed[1198],seed[3094],seed[1623],seed[1936],seed[483],seed[2075],seed[924],seed[1604],seed[3373],seed[1511],seed[2623],seed[468],seed[122],seed[1336],seed[1849],seed[4017],seed[3635],seed[456],seed[3939],seed[657],seed[3450],seed[754],seed[1894],seed[2547],seed[2792],seed[1513],seed[931],seed[1212],seed[2716],seed[2140],seed[3334],seed[3311],seed[3142],seed[2941],seed[1408],seed[3115],seed[1359],seed[672],seed[4006],seed[969],seed[279],seed[2131],seed[368],seed[1030],seed[156],seed[1628],seed[1092],seed[718],seed[3781],seed[2712],seed[2198],seed[1975],seed[262],seed[1584],seed[1761],seed[768],seed[806],seed[1892],seed[1174],seed[296],seed[1855],seed[823],seed[2927],seed[3974],seed[3436],seed[1416],seed[3993],seed[608],seed[2495],seed[3560],seed[2061],seed[3145],seed[1703],seed[2582],seed[3626],seed[1109],seed[1825],seed[2666],seed[511],seed[2281],seed[1318],seed[3850],seed[580],seed[3494],seed[3975],seed[762],seed[2887],seed[2379],seed[349],seed[106],seed[2489],seed[1521],seed[495],seed[1345],seed[3407],seed[2074],seed[778],seed[4084],seed[1167],seed[4021],seed[25],seed[1929],seed[3606],seed[3267],seed[1842],seed[564],seed[2678],seed[1564],seed[2086],seed[1870],seed[2796],seed[3364],seed[403],seed[151],seed[1726],seed[1767],seed[3394],seed[507],seed[2960],seed[1685],seed[3573],seed[1096],seed[572],seed[2451],seed[1288],seed[2209],seed[3623],seed[1962],seed[3672],seed[3228],seed[3400],seed[1832],seed[71],seed[1984],seed[324],seed[376],seed[1555],seed[3211],seed[1916],seed[1378],seed[1215],seed[234],seed[835],seed[881],seed[1042],seed[4024],seed[3237],seed[367],seed[189],seed[3163],seed[2565],seed[1502],seed[3461],seed[967],seed[137],seed[848],seed[1310],seed[2896],seed[282],seed[1873],seed[3454],seed[1989],seed[675],seed[1029],seed[571],seed[496],seed[2087],seed[482],seed[1883],seed[3717],seed[3963],seed[1142],seed[1293],seed[3528],seed[2598],seed[118],seed[1123],seed[3934],seed[742],seed[3504],seed[3133],seed[1561],seed[770],seed[1155],seed[880],seed[2311],seed[2357],seed[1931],seed[4026],seed[3527],seed[1454],seed[700],seed[1180],seed[2426],seed[2781],seed[3406],seed[3815],seed[2241],seed[1341],seed[3162],seed[1675],seed[248],seed[1444],seed[2245],seed[173],seed[170],seed[3701],seed[1247],seed[3665]}; 
//        seed7 <= {seed[426],seed[966],seed[208],seed[2963],seed[2634],seed[283],seed[4017],seed[1315],seed[2560],seed[2387],seed[1724],seed[2509],seed[927],seed[2575],seed[424],seed[2017],seed[1569],seed[3710],seed[1169],seed[2591],seed[2481],seed[1404],seed[874],seed[1491],seed[3883],seed[3967],seed[1599],seed[679],seed[676],seed[1063],seed[2138],seed[2864],seed[2825],seed[2763],seed[3460],seed[2818],seed[1791],seed[13],seed[1196],seed[1111],seed[568],seed[2292],seed[3994],seed[3351],seed[3343],seed[3073],seed[2320],seed[3765],seed[524],seed[3299],seed[3920],seed[2194],seed[1575],seed[3794],seed[1845],seed[2746],seed[3464],seed[3956],seed[3891],seed[1197],seed[2659],seed[2188],seed[1737],seed[2052],seed[1090],seed[1149],seed[2689],seed[652],seed[3328],seed[664],seed[900],seed[3595],seed[1366],seed[3761],seed[3402],seed[429],seed[2175],seed[2394],seed[445],seed[971],seed[1820],seed[736],seed[1098],seed[267],seed[1920],seed[2047],seed[3066],seed[1867],seed[3138],seed[2807],seed[1013],seed[626],seed[476],seed[2432],seed[249],seed[2754],seed[266],seed[3750],seed[151],seed[10],seed[2350],seed[852],seed[3265],seed[388],seed[1973],seed[3881],seed[2772],seed[1461],seed[2023],seed[3076],seed[3263],seed[2495],seed[841],seed[4012],seed[731],seed[138],seed[1236],seed[2987],seed[2336],seed[115],seed[3720],seed[1592],seed[4055],seed[491],seed[313],seed[1322],seed[125],seed[1529],seed[1837],seed[1226],seed[2006],seed[896],seed[2204],seed[372],seed[2829],seed[1494],seed[1789],seed[1877],seed[32],seed[1344],seed[1262],seed[1911],seed[674],seed[3626],seed[435],seed[2528],seed[2161],seed[97],seed[1495],seed[2660],seed[2348],seed[1849],seed[605],seed[3900],seed[3354],seed[3875],seed[997],seed[1385],seed[2847],seed[958],seed[1759],seed[3215],seed[2039],seed[3080],seed[2265],seed[2544],seed[906],seed[3929],seed[908],seed[62],seed[3614],seed[215],seed[2290],seed[4090],seed[2703],seed[3711],seed[3256],seed[164],seed[2679],seed[3851],seed[784],seed[411],seed[2323],seed[507],seed[1654],seed[3936],seed[3529],seed[3544],seed[3637],seed[490],seed[30],seed[2525],seed[837],seed[2124],seed[3541],seed[3699],seed[806],seed[485],seed[1132],seed[3515],seed[1878],seed[1829],seed[4025],seed[329],seed[193],seed[47],seed[203],seed[833],seed[1183],seed[348],seed[3973],seed[2142],seed[3644],seed[2295],seed[1122],seed[2782],seed[3556],seed[2379],seed[452],seed[1295],seed[1524],seed[1434],seed[2501],seed[1472],seed[1025],seed[3426],seed[600],seed[2063],seed[3240],seed[1508],seed[101],seed[1754],seed[2428],seed[2210],seed[1287],seed[3560],seed[1847],seed[1413],seed[393],seed[2885],seed[750],seed[2189],seed[3921],seed[2106],seed[1931],seed[3923],seed[2723],seed[3659],seed[3741],seed[3376],seed[3201],seed[46],seed[3686],seed[179],seed[1022],seed[1717],seed[111],seed[1251],seed[1283],seed[3648],seed[1039],seed[3363],seed[4045],seed[1813],seed[3123],seed[120],seed[683],seed[950],seed[2135],seed[2258],seed[2768],seed[3456],seed[1065],seed[812],seed[3119],seed[486],seed[1840],seed[1305],seed[2624],seed[3554],seed[1555],seed[1081],seed[3919],seed[3386],seed[102],seed[2317],seed[1735],seed[946],seed[2195],seed[409],seed[1456],seed[1546],seed[2452],seed[3745],seed[2122],seed[3910],seed[2959],seed[1469],seed[4086],seed[77],seed[2683],seed[930],seed[3840],seed[471],seed[3014],seed[2526],seed[22],seed[3521],seed[543],seed[3346],seed[3389],seed[1856],seed[1425],seed[1630],seed[140],seed[1726],seed[2310],seed[15],seed[2633],seed[3278],seed[630],seed[2981],seed[1255],seed[3597],seed[487],seed[3121],seed[2519],seed[2248],seed[1821],seed[980],seed[1916],seed[2127],seed[1927],seed[880],seed[168],seed[1693],seed[3410],seed[1384],seed[1954],seed[2021],seed[3028],seed[295],seed[2173],seed[1695],seed[1487],seed[494],seed[3372],seed[2845],seed[1997],seed[1447],seed[2190],seed[621],seed[3530],seed[1083],seed[1522],seed[1317],seed[924],seed[1518],seed[1310],seed[3142],seed[1679],seed[2249],seed[1898],seed[2802],seed[994],seed[234],seed[2433],seed[2618],seed[2539],seed[3668],seed[480],seed[3161],seed[1184],seed[3196],seed[1962],seed[3200],seed[1077],seed[3718],seed[2655],seed[3519],seed[73],seed[823],seed[2030],seed[3436],seed[3226],seed[536],seed[2028],seed[1311],seed[3636],seed[2706],seed[3949],seed[1551],seed[2270],seed[1961],seed[1335],seed[2380],seed[3183],seed[3455],seed[1258],seed[3144],seed[3168],seed[538],seed[3630],seed[3939],seed[3139],seed[3812],seed[1643],seed[2642],seed[2684],seed[1797],seed[3645],seed[2974],seed[1527],seed[3433],seed[3622],seed[651],seed[3173],seed[3228],seed[1026],seed[3442],seed[2403],seed[1362],seed[697],seed[3513],seed[2695],seed[2606],seed[2532],seed[1772],seed[3380],seed[1430],seed[12],seed[1966],seed[391],seed[3242],seed[3109],seed[2546],seed[1218],seed[1652],seed[2923],seed[1059],seed[1783],seed[37],seed[855],seed[527],seed[2902],seed[3866],seed[1155],seed[2469],seed[2031],seed[3983],seed[3149],seed[1386],seed[55],seed[2739],seed[1429],seed[2445],seed[3182],seed[1681],seed[2038],seed[1608],seed[2326],seed[1268],seed[3740],seed[2529],seed[1440],seed[776],seed[2637],seed[1248],seed[1725],seed[444],seed[3486],seed[159],seed[2698],seed[3928],seed[99],seed[1102],seed[1347],seed[3469],seed[3682],seed[1156],seed[1137],seed[1649],seed[3806],seed[1906],seed[4040],seed[2792],seed[2785],seed[1894],seed[2652],seed[3036],seed[3448],seed[3214],seed[3322],seed[2410],seed[814],seed[3338],seed[572],seed[3514],seed[71],seed[2113],seed[2430],seed[3435],seed[2828],seed[3533],seed[3255],seed[2111],seed[1776],seed[1399],seed[2202],seed[1841],seed[1061],seed[2280],seed[2774],seed[1596],seed[3086],seed[2992],seed[2570],seed[2827],seed[3826],seed[1383],seed[3972],seed[3814],seed[1237],seed[525],seed[3795],seed[1094],seed[3859],seed[314],seed[3192],seed[395],seed[530],seed[1744],seed[457],seed[364],seed[2055],seed[3285],seed[3395],seed[1235],seed[1660],seed[1123],seed[1722],seed[518],seed[3027],seed[170],seed[3450],seed[3083],seed[3445],seed[2125],seed[539],seed[341],seed[1870],seed[3500],seed[3403],seed[1680],seed[3416],seed[685],seed[3393],seed[1353],seed[1133],seed[1541],seed[2443],seed[3154],seed[1192],seed[2256],seed[3269],seed[2910],seed[2567],seed[427],seed[540],seed[1532],seed[2158],seed[2631],seed[890],seed[2592],seed[3661],seed[109],seed[942],seed[1479],seed[3052],seed[2473],seed[3522],seed[2468],seed[4093],seed[1459],seed[2770],seed[2565],seed[469],seed[4041],seed[2645],seed[260],seed[578],seed[66],seed[520],seed[1764],seed[2097],seed[1613],seed[3894],seed[337],seed[3205],seed[3749],seed[628],seed[1395],seed[3222],seed[1409],seed[3680],seed[2340],seed[3986],seed[243],seed[1466],seed[2696],seed[3494],seed[746],seed[1571],seed[1364],seed[2518],seed[2643],seed[378],seed[1401],seed[1667],seed[248],seed[2036],seed[1936],seed[2331],seed[2906],seed[2967],seed[2755],seed[2131],seed[3915],seed[1675],seed[2646],seed[1535],seed[1620],seed[2605],seed[3877],seed[2527],seed[3594],seed[478],seed[3407],seed[1993],seed[1164],seed[484],seed[380],seed[3753],seed[1828],seed[1768],seed[2579],seed[1504],seed[3047],seed[186],seed[1301],seed[3400],seed[2721],seed[563],seed[277],seed[887],seed[1860],seed[1642],seed[3227],seed[3160],seed[1588],seed[1818],seed[4032],seed[3760],seed[3441],seed[1880],seed[528],seed[1943],seed[1458],seed[3751],seed[3702],seed[1067],seed[415],seed[300],seed[2581],seed[2733],seed[2308],seed[1046],seed[3860],seed[466],seed[3114],seed[3598],seed[4023],seed[3945],seed[725],seed[1690],seed[973],seed[1050],seed[2979],seed[502],seed[3352],seed[3308],seed[253],seed[2658],seed[3037],seed[2688],seed[1068],seed[142],seed[3724],seed[3462],seed[133],seed[2497],seed[2731],seed[274],seed[3176],seed[1610],seed[270],seed[392],seed[2935],seed[1702],seed[112],seed[307],seed[1689],seed[2095],seed[1002],seed[1538],seed[1436],seed[156],seed[1810],seed[1157],seed[501],seed[2399],seed[1648],seed[3839],seed[3804],seed[35],seed[1092],seed[554],seed[3310],seed[483],seed[2298],seed[3952],seed[282],seed[3219],seed[331],seed[1908],seed[2730],seed[1583],seed[2005],seed[2788],seed[3049],seed[2145],seed[1753],seed[2100],seed[2986],seed[702],seed[2422],seed[3174],seed[2949],seed[3339],seed[2446],seed[163],seed[3298],seed[2262],seed[1874],seed[3980],seed[3022],seed[3108],seed[2781],seed[1600],seed[3854],seed[757],seed[2743],seed[2342],seed[780],seed[799],seed[1517],seed[4036],seed[926],seed[1482],seed[2933],seed[3563],seed[2182],seed[94],seed[2232],seed[1291],seed[3399],seed[2285],seed[1126],seed[872],seed[2366],seed[1162],seed[1452],seed[824],seed[1240],seed[2580],seed[1379],seed[787],seed[3535],seed[1206],seed[3373],seed[732],seed[3141],seed[1020],seed[1394],seed[3933],seed[1543],seed[3099],seed[933],seed[437],seed[3715],seed[3209],seed[1503],seed[3421],seed[303],seed[3922],seed[2835],seed[3650],seed[3788],seed[386],seed[3490],seed[3082],seed[2374],seed[1565],seed[3743],seed[2663],seed[2426],seed[2598],seed[3165],seed[3414],seed[2913],seed[3552],seed[3549],seed[2983],seed[2396],seed[1983],seed[3542],seed[3102],seed[188],seed[703],seed[717],seed[3427],seed[2457],seed[2459],seed[2700],seed[2136],seed[2744],seed[1055],seed[2453],seed[1998],seed[1418],seed[754],seed[3882],seed[2415],seed[2921],seed[3360],seed[2196],seed[643],seed[2238],seed[822],seed[959],seed[506],seed[438],seed[398],seed[2582],seed[2942],seed[3613],seed[1245],seed[1047],seed[3725],seed[2177],seed[1881],seed[1585],seed[3434],seed[3065],seed[2617],seed[1741],seed[3938],seed[2968],seed[20],seed[920],seed[1801],seed[2498],seed[4072],seed[2657],seed[2263],seed[2635],seed[3005],seed[892],seed[1963],seed[27],seed[4092],seed[516],seed[4013],seed[3169],seed[870],seed[3512],seed[2051],seed[2105],seed[2042],seed[1770],seed[192],seed[1542],seed[2397],seed[1559],seed[421],seed[58],seed[155],seed[3619],seed[2786],seed[2681],seed[2409],seed[3714],seed[219],seed[1172],seed[1121],seed[726],seed[339],seed[2960],seed[919],seed[1557],seed[3217],seed[3772],seed[1918],seed[3832],seed[646],seed[1016],seed[495],seed[982],seed[3491],seed[2260],seed[3392],seed[281],seed[3897],seed[1774],seed[1639],seed[3015],seed[3026],seed[2035],seed[2472],seed[3639],seed[1191],seed[2096],seed[577],seed[217],seed[3446],seed[2085],seed[2784],seed[1520],seed[616],seed[1799],seed[4000],seed[594],seed[1933],seed[1321],seed[2789],seed[2661],seed[448],seed[2545],seed[406],seed[3962],seed[3115],seed[1314],seed[2806],seed[2227],seed[3470],seed[3889],seed[3858],seed[2419],seed[898],seed[2141],seed[1788],seed[1892],seed[738],seed[3155],seed[2412],seed[636],seed[2651],seed[3243],seed[4043],seed[2517],seed[2090],seed[475],seed[1145],seed[917],seed[3793],seed[132],seed[3210],seed[871],seed[709],seed[2286],seed[1477],seed[1851],seed[3323],seed[1045],seed[1579],seed[3762],seed[3572],seed[3106],seed[2938],seed[1723],seed[3687],seed[2269],seed[1666],seed[645],seed[921],seed[1130],seed[3841],seed[195],seed[3095],seed[2275],seed[1578],seed[916],seed[3273],seed[2456],seed[1282],seed[3231],seed[3538],seed[2172],seed[95],seed[1342],seed[663],seed[3701],seed[410],seed[3719],seed[1330],seed[23],seed[1804],seed[811],seed[2574],seed[24],seed[2078],seed[3623],seed[2398],seed[2200],seed[653],seed[739],seed[2296],seed[1814],seed[1064],seed[3211],seed[1512],seed[701],seed[574],seed[1727],seed[113],seed[3990],seed[1400],seed[2793],seed[3982],seed[1817],seed[2108],seed[2951],seed[1439],seed[611],seed[2958],seed[3040],seed[2846],seed[867],seed[2022],seed[1378],seed[3700],seed[1739],seed[3698],seed[2471],seed[3634],seed[1533],seed[2282],seed[239],seed[1805],seed[878],seed[1471],seed[3961],seed[79],seed[2447],seed[593],seed[3705],seed[3953],seed[786],seed[2058],seed[3043],seed[2500],seed[3301],seed[3483],seed[2945],seed[2837],seed[1076],seed[2926],seed[1703],seed[316],seed[3848],seed[3580],seed[3162],seed[497],seed[2102],seed[770],seed[2319],seed[1377],seed[4037],seed[935],seed[1891],seed[265],seed[748],seed[1595],seed[3979],seed[2600],seed[756],seed[3820],seed[3046],seed[1001],seed[1843],seed[2822],seed[474],seed[1144],seed[4046],seed[3194],seed[3935],seed[623],seed[2234],seed[3093],seed[2478],seed[3291],seed[758],seed[2508],seed[1950],seed[4010],seed[2880],seed[1956],seed[52],seed[126],seed[2594],seed[141],seed[1343],seed[3452],seed[913],seed[836],seed[2899],seed[1324],seed[1165],seed[2888],seed[3768],seed[1370],seed[1298],seed[714],seed[4047],seed[1607],seed[3781],seed[981],seed[3058],seed[144],seed[199],seed[2333],seed[1771],seed[1244],seed[2450],seed[3311],seed[1574],seed[2008],seed[2347],seed[3666],seed[4027],seed[2477],seed[1286],seed[3960],seed[2084],seed[3258],seed[2114],seed[3304],seed[678],seed[3557],seed[2692],seed[695],seed[3607],seed[1826],seed[74],seed[2479],seed[2424],seed[2831],seed[2881],seed[433],seed[762],seed[2462],seed[1492],seed[1358],seed[1219],seed[268],seed[3612],seed[706],seed[418],seed[666],seed[2535],seed[114],seed[42],seed[147],seed[2046],seed[3853],seed[1116],seed[3608],seed[581],seed[1671],seed[3419],seed[569],seed[1369],seed[2146],seed[3592],seed[809],seed[216],seed[84],seed[1706],seed[988],seed[661],seed[2709],seed[1732],seed[3364],seed[2233],seed[1832],seed[3268],seed[3034],seed[2386],seed[3396],seed[365],seed[482],seed[1808],seed[3321],seed[583],seed[3097],seed[3477],seed[3502],seed[1457],seed[2395],seed[2],seed[152],seed[1309],seed[1905],seed[2454],seed[1698],seed[1035],seed[1],seed[190],seed[3569],seed[3807],seed[3199],seed[123],seed[3113],seed[2738],seed[202],seed[1118],seed[740],seed[3011],seed[2607],seed[654],seed[672],seed[3653],seed[1320],seed[1778],seed[241],seed[3633],seed[269],seed[1391],seed[1177],seed[2150],seed[470],seed[3277],seed[3378],seed[3823],seed[1949],seed[3849],seed[1955],seed[1563],seed[2727],seed[3312],seed[4071],seed[3754],seed[515],seed[2621],seed[2713],seed[2602],seed[1186],seed[2932],seed[582],seed[254],seed[2593],seed[2373],seed[720],seed[368],seed[2995],seed[3792],seed[4061],seed[3362],seed[1769],seed[2777],seed[496],seed[1684],seed[3548],seed[246],seed[1146],seed[3847],seed[1034],seed[2101],seed[1044],seed[3577],seed[1968],seed[4011],seed[1496],seed[2434],seed[3406],seed[1568],seed[2230],seed[3361],seed[259],seed[845],seed[634],seed[1940],seed[3695],seed[1308],seed[1069],seed[3135],seed[3356],seed[3536],seed[3404],seed[1719],seed[512],seed[257],seed[2192],seed[1700],seed[827],seed[2128],seed[2514],seed[3170],seed[3912],seed[3803],seed[354],seed[1141],seed[1152],seed[3420],seed[3673],seed[1110],seed[1790],seed[320],seed[3934],seed[214],seed[3041],seed[455],seed[1470],seed[3175],seed[641],seed[4015],seed[3503],seed[2247],seed[2293],seed[2082],seed[3787],seed[3487],seed[1926],seed[627],seed[2550],seed[472],seed[3329],seed[1887],seed[1590],seed[2440],seed[764],seed[1674],seed[3726],seed[2390],seed[76],seed[3625],seed[2511],seed[2823],seed[2089],seed[2564],seed[662],seed[3677],seed[2799],seed[831],seed[1350],seed[2666],seed[440],seed[135],seed[3831],seed[603],seed[608],seed[1668],seed[2538],seed[2429],seed[396],seed[2862],seed[3545],seed[2437],seed[93],seed[2253],seed[2917],seed[3507],seed[3439],seed[498],seed[1825],seed[3326],seed[3437],seed[1985],seed[2276],seed[1539],seed[3068],seed[3766],seed[3694],seed[1312],seed[1748],seed[1276],seed[1673],seed[772],seed[1420],seed[1964],seed[2029],seed[41],seed[2798],seed[3266],seed[2155],seed[119],seed[2894],seed[86],seed[304],seed[1904],seed[928],seed[2766],seed[3829],seed[1209],seed[3375],seed[960],seed[4054],seed[3481],seed[2458],seed[1979],seed[1486],seed[3588],seed[3821],seed[2185],seed[2537],seed[2726],seed[3898],seed[733],seed[1082],seed[2569],seed[1709],seed[925],seed[2874],seed[1003],seed[1972],seed[4035],seed[1793],seed[2649],seed[160],seed[103],seed[751],seed[800],seed[1593],seed[915],seed[3458],seed[2436],seed[2869],seed[3193],seed[3879],seed[2838],seed[2092],seed[918],seed[798],seed[3413],seed[951],seed[3863],seed[1975],seed[2417],seed[3264],seed[3045],seed[2499],seed[3624],seed[937],seed[2166],seed[3995],seed[3353],seed[3977],seed[251],seed[346],seed[2118],seed[3746],seed[620],seed[143],seed[2853],seed[3857],seed[2281],seed[127],seed[1037],seed[436],seed[2775],seed[2066],seed[344],seed[1502],seed[3901],seed[2217],seed[1267],seed[2669],seed[366],seed[897],seed[773],seed[2184],seed[2201],seed[2083],seed[3314],seed[1758],seed[3683],seed[3350],seed[1101],seed[3621],seed[26],seed[1526],seed[629],seed[1848],seed[3418],seed[905],seed[1659],seed[1682],seed[2912],seed[2887],seed[399],seed[3246],seed[3916],seed[3524],seed[2769],seed[3275],seed[493],seed[1318],seed[211],seed[1921],seed[3833],seed[2485],seed[213],seed[3496],seed[1188],seed[184],seed[2384],seed[3984],seed[3369],seed[4074],seed[1506],seed[2856],seed[139],seed[461],seed[3657],seed[2064],seed[308],seed[3236],seed[2000],seed[1151],seed[2555],seed[2937],seed[3180],seed[3941],seed[4018],seed[2925],seed[899],seed[1437],seed[1937],seed[3330],seed[680],seed[2294],seed[2024],seed[1902],seed[3454],seed[1000],seed[2616],seed[88],seed[2918],seed[1010],seed[2408],seed[585],seed[3651],seed[335],seed[3381],seed[1767],seed[804],seed[2324],seed[2246],seed[2274],seed[4064],seed[3056],seed[7],seed[1987],seed[2601],seed[3501],seed[3048],seed[2353],seed[1021],seed[3629],seed[3780],seed[1017],seed[4049],seed[2438],seed[499],seed[1977],seed[376],seed[3670],seed[3850],seed[3737],seed[2747],seed[2231],seed[3313],seed[408],seed[1428],seed[1269],seed[1228],seed[3493],seed[2251],seed[2257],seed[1031],seed[3129],seed[2715],seed[1323],seed[2174],seed[3830],seed[173],seed[3796],seed[1519],seed[3061],seed[1265],seed[1839],seed[730],seed[3163],seed[1270],seed[1773],seed[1895],seed[774],seed[2985],seed[2996],seed[4059],seed[271],seed[3927],seed[984],seed[673],seed[2205],seed[1550],seed[1410],seed[468],seed[224],seed[2245],seed[1942],seed[1896],seed[1525],seed[18],seed[3408],seed[955],seed[2543],seed[3985],seed[2159],seed[1742],seed[289],seed[2559],seed[548],seed[2207],seed[785],seed[579],seed[149],seed[3096],seed[1088],seed[2439],seed[3895],seed[968],seed[508],seed[521],seed[2641],seed[1302],seed[2914],seed[3571],seed[3904],seed[3835],seed[2377],seed[3307],seed[1230],seed[1463],seed[3837],seed[3184],seed[3540],seed[3239],seed[1944],seed[503],seed[1441],seed[2833],seed[3606],seed[1147],seed[2520],seed[3125],seed[1432],seed[3260],seed[204],seed[404],seed[1019],seed[2615],seed[1161],seed[2638],seed[1299],seed[3179],seed[299],seed[4038],seed[778],seed[1349],seed[1280],seed[532],seed[4044],seed[1644],seed[264],seed[1416],seed[2026],seed[3654],seed[1782],seed[3968],seed[323],seed[719],seed[82],seed[2198],seed[969],seed[877],seed[207],seed[1934],seed[1930],seed[221],seed[2832],seed[2751],seed[1627],seed[711],seed[3691],seed[4006],seed[340],seed[1890],seed[1665],seed[3116],seed[1140],seed[1057],seed[2972],seed[2506],seed[158],seed[4091],seed[178],seed[2778],seed[2370],seed[2123],seed[1755],seed[2240],seed[3635],seed[1548],seed[3476],seed[4057],seed[614],seed[2599],seed[0],seed[2924],seed[2402],seed[3131],seed[453],seed[130],seed[2783],seed[2327],seed[660],seed[2305],seed[2512],seed[328],seed[302],seed[1204],seed[1852],seed[1919],seed[3672],seed[136],seed[2557],seed[2041],seed[3267],seed[2465],seed[306],seed[745],seed[1408],seed[50],seed[2991],seed[3417],seed[1928],seed[2164],seed[1868],seed[1691],seed[941],seed[3128],seed[2842],seed[3627],seed[1711],seed[1696],seed[2699],seed[3012],seed[454],seed[2705],seed[2801],seed[4069],seed[1053],seed[4030],seed[866],seed[1327],seed[1996],seed[1345],seed[2109],seed[1093],seed[4065],seed[2416],seed[1078],seed[2153],seed[3603],seed[183],seed[4066],seed[2455],seed[1728],seed[1040],seed[3689],seed[353],seed[1091],seed[3252],seed[834],seed[90],seed[3996],seed[954],seed[1952],seed[2040],seed[2065],seed[3038],seed[965],seed[3358],seed[3855],seed[3728],seed[847],seed[3827],seed[696],seed[983],seed[1337],seed[808],seed[3447],seed[1483],seed[1333],seed[3534],seed[1313],seed[3091],seed[2757],seed[2736],seed[2015],seed[3300],seed[617],seed[670],seed[129],seed[3674],seed[3394],seed[3523],seed[1749],seed[389],seed[294],seed[1213],seed[1765],seed[2886],seed[1641],seed[2664],seed[401],seed[881],seed[3468],seed[850],seed[1806],seed[1917],seed[715],seed[3148],seed[3575],seed[2405],seed[2989],seed[458],seed[3218],seed[3000],seed[952],seed[263],seed[551],seed[49],seed[1227],seed[3744],seed[360],seed[637],seed[1498],seed[4014],seed[2662],seed[2139],seed[2909],seed[1351],seed[2577],seed[1406],seed[3002],seed[2898],seed[2704],seed[1969],seed[2361],seed[3690],seed[2915],seed[3325],seed[1072],seed[1203],seed[456],seed[1398],seed[59],seed[3574],seed[3401],seed[324],seed[2488],seed[598],seed[3786],seed[2507],seed[1234],seed[318],seed[633],seed[665],seed[595],seed[325],seed[379],seed[1951],seed[2316],seed[2104],seed[2053],seed[1734],seed[3620],seed[33],seed[3459],seed[1297],seed[3824],seed[349],seed[3931],seed[622],seed[3669],seed[1655],seed[3319],seed[2197],seed[1217],seed[1631],seed[1014],seed[909],seed[1882],seed[2761],seed[3596],seed[4068],seed[167],seed[2750],seed[3112],seed[2191],seed[604],seed[2558],seed[131],seed[319],seed[3771],seed[2977],seed[3188],seed[280],seed[1611],seed[3678],seed[1511],seed[2572],seed[3225],seed[1307],seed[4026],seed[3411],seed[3911],seed[1705],seed[3940],seed[953],seed[1553],seed[2648],seed[1290],seed[227],seed[2335],seed[489],seed[3963],seed[3294],seed[137],seed[2855],seed[89],seed[1685],seed[244],seed[3092],seed[3553],seed[1999],seed[2562],seed[1859],seed[1154],seed[3449],seed[1490],seed[3805],seed[276],seed[220],seed[1075],seed[510],seed[500],seed[2813],seed[3136],seed[1087],seed[2144],seed[3247],seed[1277],seed[1259],seed[2300],seed[2115],seed[3782],seed[1249],seed[707],seed[1124],seed[2765],seed[3430],seed[2267],seed[2608],seed[3685],seed[2866],seed[1194],seed[613],seed[181],seed[3006],seed[2208],seed[326],seed[4052],seed[3903],seed[2423],seed[1266],seed[2759],seed[3366],seed[2032],seed[2536],seed[2264],seed[355],seed[1853],seed[3282],seed[995],seed[361],seed[2461],seed[1854],seed[296],seed[1816],seed[1449],seed[1085],seed[2140],seed[4020],seed[3584],seed[148],seed[1547],seed[1971],seed[1581],seed[2919],seed[1285],seed[3074],seed[2463],seed[460],seed[549],seed[1095],seed[1617],seed[3886],seed[1125],seed[3089],seed[434],seed[1857],seed[2676],seed[2199],seed[1105],seed[1360],seed[1444],seed[1530],seed[1205],seed[1795],seed[1626],seed[3551],seed[4088],seed[3079],seed[3861],seed[2072],seed[3758],seed[397],seed[1923],seed[3717],seed[3951],seed[1293],seed[2425],seed[2007],seed[3457],seed[1056],seed[2540],seed[1893],seed[638],seed[3133],seed[1422],seed[3050],seed[2805],seed[105],seed[2012],seed[943],seed[655],seed[843],seed[1241],seed[708],seed[2711],seed[1243],seed[1913],seed[3713],seed[3943],seed[1558],seed[1182],seed[2844],seed[553],seed[816],seed[1780],seed[3932],seed[2762],seed[2929],seed[3062],seed[3601],seed[3706],seed[3561],seed[2057],seed[2836],seed[226],seed[1621],seed[237],seed[2219],seed[2928],seed[2206],seed[3018],seed[2753],seed[2119],seed[904],seed[3884],seed[1319],seed[3398],seed[2742],seed[741],seed[3819],seed[2796],seed[3518],seed[3759],seed[1138],seed[3974],seed[2586],seed[3573],seed[3384],seed[2722],seed[1763],seed[2381],seed[407],seed[1250],seed[2302],seed[25],seed[1339],seed[1256],seed[1338],seed[1619],seed[3024],seed[3785],seed[2841],seed[2604],seed[1622],seed[54],seed[3206],seed[3259],seed[911],seed[2020],seed[1827],seed[3517],seed[1128],seed[402],seed[367],seed[687],seed[934],seed[2952],seed[1946],seed[3289],seed[3516],seed[3585],seed[1396],seed[2080],seed[2566],seed[2213],seed[2087],seed[3021],seed[2901],seed[2002],seed[3838],seed[1272],seed[3492],seed[768],seed[3320],seed[882],seed[2800],seed[1594],seed[1907],seed[3071],seed[3122],seed[1214],seed[990],seed[3388],seed[3118],seed[1865],seed[3693],seed[3475],seed[3808],seed[2611],seed[3482],seed[1986],seed[3582],seed[1640],seed[3371],seed[3937],seed[3315],seed[4083],seed[3647],seed[667],seed[876],seed[315],seed[2266],seed[1390],seed[2033],seed[755],seed[2625],seed[2130],seed[122],seed[1591],seed[180],seed[3212],seed[2309],seed[3060],seed[596],seed[1454],seed[1570],seed[2549],seed[3905],seed[1080],seed[3004],seed[145],seed[3473],seed[209],seed[2225],seed[3907],seed[403],seed[3716],seed[1796],seed[2418],seed[2167],seed[2341],seed[2045],seed[3656],seed[828],seed[229],seed[1721],seed[2834],seed[795],seed[3667],seed[428],seed[4004],seed[698],seed[2067],seed[75],seed[2226],seed[169],seed[100],seed[3409],seed[3337],seed[1150],seed[1348],seed[3570],seed[2851],seed[519],seed[3727],seed[1381],seed[609],seed[3357],seed[1274],seed[1509],seed[1208],seed[1402],seed[3997],seed[431],seed[657],seed[3098],seed[2328],seed[2810],seed[825],seed[631],seed[118],seed[2103],seed[87],seed[2815],seed[2363],seed[1794],seed[2411],seed[2980],seed[1024],seed[2487],seed[3971],seed[1015],seed[2668],seed[2767],seed[1008],seed[1629],seed[2362],seed[1216],seed[979],seed[2486],seed[597],seed[3547],seed[844],seed[4048],seed[1393],seed[2148],seed[505],seed[1670],seed[936],seed[245],seed[2367],seed[3164],seed[2356],seed[2571],seed[3334],seed[1117],seed[3213],seed[53],seed[2365],seed[3077],seed[3488],seed[2489],seed[647],seed[298],seed[2156],seed[272],seed[3262],seed[3423],seed[3377],seed[2171],seed[1468],seed[3137],seed[3132],seed[2587],seed[1423],seed[3472],seed[1787],seed[1683],seed[2165],seed[345],seed[2371],seed[1676],seed[1582],seed[3117],seed[3834],seed[327],seed[382],seed[2982],seed[3987],seed[3140],seed[2719],seed[3237],seed[1612],seed[417],seed[2680],seed[2435],seed[39],seed[3739],seed[4078],seed[3942],seed[1751],seed[3153],seed[691],seed[846],seed[964],seed[284],seed[2953],seed[1862],seed[2523],seed[200],seed[902],seed[146],seed[2843],seed[3784],seed[601],seed[198],seed[1537],seed[2081],seed[888],seed[1359],seed[526],seed[2242],seed[3899],seed[879],seed[564],seed[818],seed[2858],seed[2152],seed[3280],seed[252],seed[1939],seed[1252],seed[1688],seed[2406],seed[2650],seed[1033],seed[618],seed[3611],seed[2884],seed[1633],seed[2734],seed[4005],seed[36],seed[2277],seed[1103],seed[2613],seed[1435],seed[1442],seed[1296],seed[565],seed[2522],seed[791],seed[1325],seed[2315],seed[863],seed[3978],seed[1647],seed[2444],seed[1462],seed[369],seed[3391],seed[796],seed[793],seed[3478],seed[3800],seed[1635],seed[835],seed[976],seed[1304],seed[3511],seed[171],seed[1586],seed[2687],seed[261],seed[588],seed[3688],seed[1989],seed[1836],seed[3272],seed[523],seed[649],seed[2916],seed[174],seed[961],seed[561],seed[17],seed[3223],seed[78],seed[2821],seed[1238],seed[1136],seed[895],seed[759],seed[2712],seed[2547],seed[2623],seed[4075],seed[1179],seed[749],seed[586],seed[1699],seed[2513],seed[1131],seed[3872],seed[3589],seed[1779],seed[684],seed[560],seed[813],seed[1510],seed[1980],seed[1200],seed[3064],seed[124],seed[729],seed[177],seed[2301],seed[3425],seed[2717],seed[535],seed[3370],seed[416],seed[3506],seed[4007],seed[3017],seed[2748],seed[3202],seed[977],seed[1866],seed[688],seed[3846],seed[752],seed[154],seed[2797],seed[446],seed[3059],seed[2493],seed[2957],seed[893],seed[1375],seed[802],seed[150],seed[765],seed[3382],seed[587],seed[3809],seed[3467],seed[3432],seed[2947],seed[405],seed[2160],seed[639],seed[1176],seed[3293],seed[1809],seed[1160],seed[700],seed[1864],seed[3776],seed[1411],seed[2872],seed[1397],seed[3085],seed[2337],seed[3964],seed[2203],seed[3220],seed[1480],seed[2988],seed[2521],seed[3681],seed[840],seed[1750],seed[1222],seed[3662],seed[1861],seed[2510],seed[1833],seed[3063],seed[2737],seed[2503],seed[1900],seed[3100],seed[2391],seed[2883],seed[1300],seed[632],seed[1807],seed[2178],seed[2376],seed[3198],seed[1499],seed[2678],seed[1746],seed[1005],seed[3692],seed[3271],seed[2708],seed[4062],seed[713],seed[1048],seed[2812],seed[2393],seed[2025],seed[2218],seed[537],seed[1991],seed[3224],seed[2795],seed[2170],seed[414],seed[2466],seed[2496],seed[3887],seed[1210],seed[117],seed[1340],seed[2873],seed[1104],seed[2330],seed[3498],seed[3345],seed[1143],seed[658],seed[3822],seed[4033],seed[1071],seed[3107],seed[3738],seed[333],seed[2934],seed[1284],seed[914],seed[3281],seed[305],seed[4001],seed[3583],seed[838],seed[44],seed[2716],seed[2877],seed[1863],seed[3587],seed[2287],seed[1978],seed[656],seed[681],seed[2970],seed[1198],seed[2318],seed[210],seed[2420],seed[1855],seed[3958],seed[2349],seed[1577],seed[2237],seed[2404],seed[1038],seed[1948],seed[2427],seed[2780],seed[2414],seed[2186],seed[3365],seed[2946],seed[2378],seed[2223],seed[2329],seed[1148],seed[1485],seed[3537],seed[2961],seed[1914],seed[3642],seed[1786],seed[989],seed[1374],seed[3344],seed[1775],seed[1616],seed[3546],seed[383],seed[3124],seed[92],seed[514],seed[1701],seed[373],seed[699],seed[1412],seed[3852],seed[317],seed[3250],seed[884],seed[3504],seed[3296],seed[342],seed[807],seed[3254],seed[1231],seed[2311],seed[3185],seed[1982],seed[3248],seed[3764],seed[2034],seed[3777],seed[2840],seed[357],seed[1306],seed[425],seed[3075],seed[3126],seed[68],seed[1784],seed[1481],seed[1012],seed[2355],seed[3429],seed[3729],seed[2504],seed[1835],seed[689],seed[2074],seed[492],seed[3813],seed[3147],seed[1253],seed[2049],seed[3825],seed[2241],seed[2922],seed[3558],seed[3039],seed[3505],seed[8],seed[2235],seed[1731],seed[4094],seed[3348],seed[2773],seed[1716],seed[3324],seed[2401],seed[3618],seed[1965],seed[3244],seed[2892],seed[2860],seed[96],seed[3461],seed[3568],seed[3665],seed[753],seed[1545],seed[3238],seed[2011],seed[975],seed[3525],seed[1168],seed[419],seed[1058],seed[3908],seed[2895],seed[2261],seed[1598],seed[734],seed[3203],seed[682],seed[2876],seed[949],seed[1247],seed[3615],seed[2467],seed[377],seed[166],seed[3902],seed[3721],seed[1678],seed[1451],seed[1850],seed[2464],seed[3555],seed[1792],seed[2553],seed[1229],seed[225],seed[1041],seed[1812],seed[232],seed[3871],seed[1326],seed[932],seed[1561],seed[297],seed[1341],seed[1007],seed[3870],seed[2820],seed[2694],seed[2997],seed[1677],seed[1514],seed[2243],seed[1139],seed[550],seed[3335],seed[3485],seed[1536],seed[3390],seed[3158],seed[247],seed[2729],seed[2875],seed[1281],seed[3969],seed[939],seed[1417],seed[1988],seed[1687],seed[3207],seed[4021],seed[412],seed[1938],seed[2707],seed[288],seed[473],seed[974],seed[1084],seed[3428],seed[1450],seed[2181],seed[2573],seed[3438],seed[1257],seed[9],seed[31],seed[3867],seed[3290],seed[1329],seed[287],seed[3251],seed[826],seed[829],seed[2891],seed[944],seed[612],seed[889],seed[1884],seed[801],seed[3208],seed[1356],seed[2597],seed[602],seed[1540],seed[222],seed[2289],seed[3649],seed[1875],seed[865],seed[3991],seed[2870],seed[2480],seed[1279],seed[3181],seed[2303],seed[1263],seed[513],seed[3736],seed[3842],seed[423],seed[2852],seed[1941],seed[3906],seed[1576],seed[3696],seed[3609],seed[1883],seed[3981],seed[2673],seed[1730],seed[2516],seed[1844],seed[985],seed[2896],seed[1811],seed[2009],seed[3177],seed[2279],seed[692],seed[1185],seed[3055],seed[2760],seed[2126],seed[504],seed[967],seed[2561],seed[2069],seed[2897],seed[886],seed[3733],seed[2339],seed[3233],seed[3104],seed[3712],seed[29],seed[3463],seed[1066],seed[301],seed[2010],seed[763],seed[2848],seed[1516],seed[3397],seed[1175],seed[1135],seed[3799],seed[1163],seed[2907],seed[3874],seed[1625],seed[1521],seed[862],seed[2332],seed[3235],seed[3495],seed[3878],seed[347],seed[6],seed[2644],seed[1387],seed[63],seed[462],seed[3274],seed[2344],seed[2304],seed[2563],seed[3641],seed[3042],seed[2273],seed[978],seed[2619],seed[3815],seed[1580],seed[3292],seed[2120],seed[3646],seed[4067],seed[3489],seed[3016],seed[4009],seed[3527],seed[1294],seed[3306],seed[571],seed[2674],seed[1011],seed[1223],seed[238],seed[3697],seed[1328],seed[1967],seed[2656],seed[3888],seed[1947],seed[693],seed[1365],seed[894],seed[2849],seed[4073],seed[2050],seed[3305],seed[2505],seed[2578],seed[2596],seed[625],seed[3566],seed[2086],seed[1407],seed[1756],seed[1505],seed[3443],seed[769],seed[273],seed[2830],seed[2244],seed[191],seed[2530],seed[2839],seed[2076],seed[1995],seed[3303],seed[2059],seed[782],seed[3783],seed[3845],seed[3660],seed[710],seed[439],seed[1872],seed[3287],seed[2998],seed[3676],seed[2622],seed[992],seed[3811],seed[1166],seed[3703],seed[1464],seed[2474],seed[3959],seed[875],seed[2077],seed[2603],seed[64],seed[3671],seed[359],seed[3284],seed[2112],seed[285],seed[3288],seed[3790],seed[1260],seed[2252],seed[1858],seed[2070],seed[3031],seed[998],seed[2271],seed[3638],seed[321],seed[947],seed[3166],seed[1924],seed[3054],seed[957],seed[1707],seed[3734],seed[2117],seed[2590],seed[1632],seed[1573],seed[2941],seed[1604],seed[2654],seed[3869],seed[3105],seed[2451],seed[2180],seed[2677],seed[91],seed[1662],seed[2272],seed[48],seed[3216],seed[3032],seed[2359],seed[2375],seed[2056],seed[3893],seed[4070],seed[742],seed[2697],seed[690],seed[3509],seed[2809],seed[2460],seed[1113],seed[2944],seed[3286],seed[3159],seed[1889],seed[573],seed[57],seed[1745],seed[1932],seed[2220],seed[28],seed[2609],seed[589],seed[1424],seed[2690],seed[2037],seed[3090],seed[1115],seed[3775],seed[2048],seed[2653],seed[189],seed[3778],seed[907],seed[3270],seed[2013],seed[1556],seed[1747],seed[2610],seed[4024],seed[4058],seed[3543],seed[443],seed[1661],seed[3909],seed[1086],seed[3081],seed[744],seed[2714],seed[420],seed[1515],seed[2826],seed[1615],seed[712],seed[1193],seed[2254],seed[2640],seed[1567],seed[624],seed[3088],seed[1752],seed[590],seed[2595],seed[1692],seed[2369],seed[3331],seed[1389],seed[2808],seed[1336],seed[3652],seed[3999],seed[948],seed[1489],seed[2211],seed[2016],seed[3632],seed[1802],seed[3789],seed[387],seed[488],seed[4034],seed[34],seed[3631],seed[2556],seed[3072],seed[3828],seed[3600],seed[3617],seed[2321],seed[2133],seed[3966],seed[116],seed[1766],seed[1651],seed[21],seed[3257],seed[1669],seed[1478],seed[3843],seed[3355],seed[4016],seed[206],seed[4019],seed[3151],seed[901],seed[558],seed[3890],seed[2639],seed[3466],seed[619],seed[1376],seed[2222],seed[2728],seed[3559],seed[1030],seed[566],seed[3810],seed[2632],seed[128],seed[336],seed[2554],seed[1736],seed[3057],seed[3892],seed[1974],seed[1465],seed[1733],seed[1431],seed[727],seed[1029],seed[3013],seed[2228],seed[107],seed[1672],seed[4089],seed[2614],seed[2911],seed[4],seed[240],seed[1028],seed[233],seed[2392],seed[803],seed[1901],seed[3992],seed[517],seed[671],seed[790],seed[197],seed[1049],seed[3019],seed[1473],seed[747],seed[987],seed[1929],seed[1899],seed[533],seed[938],seed[2221],seed[559],seed[3033],seed[1623],seed[3709],seed[2268],seed[2132],seed[1710],seed[2068],seed[1953],seed[371],seed[591],seed[3143],seed[3988],seed[3748],seed[1445],seed[3276],seed[1224],seed[555],seed[467],seed[1497],seed[3586],seed[3955],seed[2857],seed[3035],seed[1242],seed[3773],seed[2954],seed[2824],seed[3742],seed[218],seed[3010],seed[2701],seed[2948],seed[1142],seed[2491],seed[922],seed[2627],seed[1114],seed[3581],seed[686],seed[134],seed[3309],seed[3924],seed[839],seed[2749],seed[1712],seed[1054],seed[2670],seed[1127],seed[3918],seed[2183],seed[1523],seed[2179],seed[2325],seed[14],seed[2382],seed[104],seed[1189],seed[669],seed[3186],seed[2740],seed[1822],seed[358],seed[3453],seed[3152],seed[2307],seed[2969],seed[3383],seed[4042],seed[3341],seed[704],seed[2879],seed[1361],seed[1448],seed[3976],seed[694],seed[2278],seed[3970],seed[3679],seed[1597],seed[1158],seed[1460],seed[310],seed[3431],seed[2551],seed[2850],seed[858],seed[394],seed[2043],seed[2389],seed[3230],seed[2667],seed[1572],seed[2388],seed[2482],seed[3003],seed[1475],seed[2920],seed[3684],seed[375],seed[2718],seed[547],seed[2685],seed[2956],seed[606],seed[1658],seed[1903],seed[4003],seed[1992],seed[3150],seed[2091],seed[2413],seed[1871],seed[1879],seed[1686],seed[1488],seed[3261],seed[2671],seed[1120],seed[1781],seed[2620],seed[2476],seed[83],seed[821],seed[2647],seed[760],seed[3479],seed[2368],seed[562],seed[1609],seed[3379],seed[1079],seed[4053],seed[1885],seed[635],seed[1371],seed[2383],seed[390],seed[1199],seed[3655],seed[2116],seed[1190],seed[2149],seed[3747],seed[1036],seed[81],seed[2098],seed[2475],seed[3767],seed[290],seed[1886],seed[72],seed[2019],seed[2939],seed[1419],seed[1443],seed[3295],seed[1346],seed[1645],seed[860],seed[1562],seed[962],seed[3008],seed[1352],seed[923],seed[3658],seed[1415],seed[1211],seed[286],seed[1264],seed[2214],seed[945],seed[1664],seed[463],seed[724],seed[3510],seed[3816],seed[3007],seed[3817],seed[3101],seed[2965],seed[3730],seed[1564],seed[1708],seed[4056],seed[2004],seed[2212],seed[309],seed[370],seed[956],seed[2283],seed[2568],seed[38],seed[1650],seed[3249],seed[3868],seed[1761],seed[1922],seed[737],seed[3593],seed[2930],seed[2284],seed[2993],seed[1382],seed[3067],seed[356],seed[1292],seed[1606],seed[1657],seed[2001],seed[869],seed[3318],seed[2364],seed[1178],seed[910],seed[1427],seed[2215],seed[3440],seed[3084],seed[2421],seed[972],seed[963],seed[2542],seed[1785],seed[1873],seed[2297],seed[2533],seed[3539],seed[2110],seed[2431],seed[3732],seed[2900],seed[3191],seed[2407],seed[3451],seed[1601],seed[777],seed[278],seed[1354],seed[1388],seed[255],seed[3023],seed[441],seed[883],seed[2863],seed[3070],seed[3770],seed[1958],seed[3221],seed[1212],seed[3774],seed[2003],seed[3779],seed[1027],seed[2752],seed[644],seed[3708],seed[820],seed[3],seed[1912],seed[2314],seed[2994],seed[2745],seed[2187],seed[4079],seed[172],seed[4076],seed[1438],seed[575],seed[1099],seed[2682],seed[3178],seed[1106],seed[2163],seed[1528],seed[1959],seed[2306],seed[1221],seed[2758],seed[3722],seed[175],seed[3332],seed[3914],seed[352],seed[931],seed[2176],seed[3550],seed[1976],seed[5],seed[1180],seed[293],seed[2490],seed[4085],seed[761],seed[3387],seed[3336],seed[374],seed[3317],seed[3565],seed[991],seed[2971],seed[797],seed[2675],seed[2062],seed[1119],seed[3359],seed[351],seed[311],seed[2027],seed[3531],seed[640],seed[929],seed[3241],seed[2484],seed[2903],seed[856],seed[3197],seed[3798],seed[1170],seed[2515],seed[2976],seed[1070],seed[3755],seed[1697],seed[1738],seed[650],seed[1009],seed[940],seed[1476],seed[873],seed[1373],seed[1004],seed[1246],seed[1876],seed[3316],seed[542],seed[1815],seed[3349],seed[842],seed[2054],seed[1614],seed[1638],seed[4008],seed[2854],seed[2966],seed[3094],seed[567],seed[43],seed[1403],seed[3499],seed[153],seed[1051],seed[2216],seed[3801],seed[3975],seed[3769],seed[552],seed[3030],seed[3465],seed[3497],seed[735],seed[1605],seed[4039],seed[2882],seed[2531],seed[3422],seed[194],seed[1042],seed[3526],seed[781],seed[3156],seed[2441],seed[2259],seed[1129],seed[1074],seed[3731],seed[3171],seed[1357],seed[851],seed[40],seed[464],seed[2904],seed[1842],seed[69],seed[2137],seed[3412],seed[2867],seed[3145],seed[2018],seed[1453],seed[1271],seed[2352],seed[2771],seed[1023],seed[3599],seed[1869],seed[3110],seed[3025],seed[2168],seed[362],seed[2732],seed[534],seed[2162],seed[2372],seed[3913],seed[1720],seed[3528],seed[1363],seed[442],seed[2779],seed[1910],seed[2483],seed[2878],seed[2470],seed[1355],seed[2552],seed[2962],seed[3297],seed[4060],seed[3604],seed[2134],seed[1159],seed[1233],seed[1646],seed[1513],seed[2343],seed[832],seed[1501],seed[1824],seed[1714],seed[3001],seed[2071],seed[767],seed[903],seed[3930],seed[2589],seed[1426],seed[2079],seed[912],seed[80],seed[3232],seed[3602],seed[3757],seed[291],seed[2583],seed[675],seed[2816],seed[1367],seed[779],seed[3675],seed[1334],seed[201],seed[2358],seed[3484],seed[2725],seed[3643],seed[1331],seed[2693],seed[1153],seed[4080],seed[250],seed[2803],seed[993],seed[1405],seed[4050],seed[3917],seed[106],seed[2794],seed[3965],seed[2313],seed[810],seed[2291],seed[3865],seed[2229],seed[1018],seed[3333],seed[1500],seed[531],seed[2494],seed[3053],seed[2044],seed[599],seed[1945],seed[2636],seed[1220],seed[576],seed[610],seed[970],seed[2905],seed[3947],seed[1994],seed[1743],seed[2819],seed[2585],seed[2859],seed[3134],seed[235],seed[3342],seed[2448],seed[343],seed[4051],seed[182],seed[2129],seed[3130],seed[864],seed[1960],seed[3993],seed[1109],seed[381],seed[1062],seed[3948],seed[479],seed[1332],seed[1507],seed[2239],seed[1800],seed[556],seed[1052],seed[2099],seed[2984],seed[70],seed[4081],seed[2107],seed[422],seed[509],seed[1207],seed[2088],seed[67],seed[60],seed[3957],seed[1587],seed[2628],seed[1421],seed[3157],seed[2990],seed[3616],seed[2868],seed[275],seed[642],seed[1534],seed[3187],seed[3567],seed[3864],seed[1990],seed[1134],seed[450],seed[1544],seed[1715],seed[3532],seed[196],seed[165],seed[11],seed[3253],seed[2385],seed[262],seed[857],seed[2940],seed[2764],seed[447],seed[1618],seed[2400],seed[1275],seed[1628],seed[848],seed[1089],seed[2691],seed[400],seed[522],seed[789],seed[3204],seed[228],seed[999],seed[1925],seed[4087],seed[1554],seed[677],seed[1602],seed[868],seed[110],seed[2710],seed[2927],seed[4022],seed[541],seed[3954],seed[2534],seed[3880],seed[1288],seed[1167],seed[854],seed[384],seed[432],seed[161],seed[3368],seed[1566],seed[1589],seed[1549],seed[545],seed[4084],seed[1372],seed[1195],seed[3245],seed[1834],seed[3229],seed[1202],seed[2502],seed[3578],seed[3424],seed[1729],seed[3876],seed[859],seed[1984],seed[3576],seed[2147],seed[1757],seed[1718],seed[788],seed[3195],seed[3103],seed[4029],seed[2865],seed[1225],seed[2255],seed[3836],seed[1560],seed[242],seed[3127],seed[794],seed[2157],seed[721],seed[986],seed[1909],seed[668],seed[3763],seed[1368],seed[1455],seed[2955],seed[1915],seed[413],seed[570],seed[465],seed[205],seed[108],seed[2312],seed[2169],seed[3146],seed[2346],seed[350],seed[2686],seed[1694],seed[511],seed[363],seed[332],seed[2014],seed[2061],seed[3707],seed[223],seed[1201],seed[3562],seed[1073],seed[230],seed[1303],seed[3340],seed[1232],seed[1107],seed[61],seed[2121],seed[891],seed[3885],seed[1278],seed[3925],seed[3009],seed[3640],seed[1713],seed[728],seed[3896],seed[121],seed[322],seed[3167],seed[3234],seed[792],seed[830],seed[1108],seed[3520],seed[236],seed[3862],seed[2814],seed[805],seed[2250],seed[2629],seed[2449],seed[722],seed[3926],seed[2576],seed[2151],seed[783],seed[176],seed[330],seed[258],seed[2790],seed[1803],seed[2908],seed[1289],seed[1187],seed[3756],seed[3590],seed[1935],seed[1762],seed[3405],seed[1096],seed[4002],seed[705],seed[2588],seed[157],seed[1760],seed[3078],seed[3374],seed[4082],seed[385],seed[3471],seed[718],seed[3591],seed[2665],seed[2338],seed[2964],seed[607],seed[430],seed[2584],seed[1174],seed[3797],seed[2073],seed[1173],seed[2999],seed[2931],seed[4095],seed[659],seed[557],seed[19],seed[1484],seed[1603],seed[3508],seed[2357],seed[592],seed[815],seed[231],seed[885],seed[2861],seed[1215],seed[3069],seed[1392],seed[580],seed[3723],seed[3844],seed[2236],seed[1634],seed[338],seed[2811],seed[1261],seed[3279],seed[2360],seed[3989],seed[2548],seed[1552],seed[2322],seed[2936],seed[3051],seed[1060],seed[477],seed[2893],seed[1798],seed[3283],seed[2060],seed[4063],seed[648],seed[861],seed[2154],seed[2817],seed[2143],seed[2943],seed[334],seed[544],seed[743],seed[1663],seed[2890],seed[3172],seed[1097],seed[1032],seed[2351],seed[853],seed[1446],seed[279],seed[1831],seed[1636],seed[817],seed[716],seed[2209],seed[1006],seed[65],seed[2354],seed[2791],seed[2787],seed[2756],seed[2094],seed[3610],seed[4028],seed[16],seed[85],seed[2889],seed[819],seed[1273],seed[1433],seed[1653],seed[3087],seed[3818],seed[849],seed[1656],seed[292],seed[3474],seed[1897],seed[2442],seed[1740],seed[1043],seed[2299],seed[459],seed[1171],seed[2776],seed[1239],seed[1414],seed[1981],seed[451],seed[56],seed[2288],seed[3189],seed[3020],seed[4077],seed[1777],seed[2075],seed[3950],seed[1474],seed[1970],seed[45],seed[2720],seed[1316],seed[3385],seed[2804],seed[775],seed[584],seed[185],seed[2224],seed[162],seed[2735],seed[3367],seed[1380],seed[3735],seed[481],seed[2871],seed[4031],seed[2702],seed[2978],seed[3302],seed[3791],seed[3579],seed[2524],seed[3663],seed[3111],seed[2334],seed[98],seed[2541],seed[2975],seed[771],seed[3664],seed[1100],seed[1584],seed[1830],seed[1823],seed[3190],seed[1957],seed[1819],seed[3347],seed[3605],seed[3873],seed[2741],seed[2612],seed[2492],seed[1704],seed[546],seed[3998],seed[1624],seed[723],seed[3029],seed[3856],seed[3944],seed[51],seed[1531],seed[766],seed[2950],seed[212],seed[187],seed[1112],seed[3444],seed[449],seed[996],seed[3802],seed[3327],seed[2093],seed[2973],seed[256],seed[1888],seed[2345],seed[3752],seed[312],seed[3946],seed[1181],seed[3480],seed[1493],seed[2724],seed[3564],seed[2672],seed[1467],seed[615],seed[3704],seed[529],seed[1637],seed[1254],seed[2193],seed[3415],seed[3044],seed[2630],seed[2626],seed[1838],seed[1846],seed[3628],seed[3120]}; 
//        seed8 <= {seed[2128],seed[2719],seed[1599],seed[3598],seed[1369],seed[1503],seed[1622],seed[241],seed[2621],seed[1680],seed[2037],seed[3670],seed[3210],seed[3434],seed[3846],seed[22],seed[3829],seed[2936],seed[2283],seed[1910],seed[1088],seed[3817],seed[462],seed[3080],seed[1689],seed[3419],seed[150],seed[1999],seed[273],seed[957],seed[3488],seed[1798],seed[1460],seed[3892],seed[1277],seed[3740],seed[2261],seed[3403],seed[2206],seed[1959],seed[255],seed[2183],seed[504],seed[3681],seed[2625],seed[2184],seed[3145],seed[1579],seed[3156],seed[3855],seed[2990],seed[2319],seed[2314],seed[2321],seed[4081],seed[3966],seed[1373],seed[1051],seed[2536],seed[2058],seed[2520],seed[989],seed[2696],seed[3352],seed[565],seed[92],seed[3591],seed[2138],seed[2063],seed[2578],seed[1748],seed[1279],seed[956],seed[60],seed[3884],seed[2948],seed[2142],seed[1254],seed[1833],seed[455],seed[2710],seed[2714],seed[2753],seed[1333],seed[1349],seed[2407],seed[1614],seed[2020],seed[1233],seed[3602],seed[2734],seed[550],seed[1451],seed[673],seed[4058],seed[1228],seed[2120],seed[1640],seed[3933],seed[2046],seed[1057],seed[3465],seed[2608],seed[2829],seed[18],seed[1371],seed[3249],seed[1558],seed[2452],seed[3706],seed[1027],seed[703],seed[1884],seed[269],seed[864],seed[2295],seed[2551],seed[3504],seed[2950],seed[441],seed[2945],seed[2332],seed[927],seed[2777],seed[2679],seed[2790],seed[928],seed[3556],seed[2723],seed[2126],seed[3848],seed[1975],seed[1453],seed[1791],seed[1545],seed[6],seed[1583],seed[171],seed[2351],seed[2820],seed[522],seed[1463],seed[1977],seed[1040],seed[3734],seed[3317],seed[2812],seed[3111],seed[1025],seed[1500],seed[373],seed[1416],seed[3195],seed[2534],seed[629],seed[606],seed[1817],seed[3801],seed[1571],seed[595],seed[2703],seed[839],seed[3028],seed[2430],seed[1075],seed[562],seed[1466],seed[3522],seed[238],seed[1816],seed[614],seed[915],seed[2403],seed[2983],seed[2417],seed[2739],seed[648],seed[110],seed[2494],seed[2080],seed[714],seed[2911],seed[2055],seed[712],seed[2047],seed[807],seed[3297],seed[3222],seed[936],seed[1178],seed[3004],seed[1395],seed[3753],seed[3112],seed[157],seed[3253],seed[1449],seed[2666],seed[1674],seed[2081],seed[878],seed[95],seed[2862],seed[1273],seed[615],seed[3225],seed[2641],seed[1157],seed[1991],seed[530],seed[2467],seed[2928],seed[2560],seed[2962],seed[2176],seed[3068],seed[676],seed[747],seed[3362],seed[474],seed[3940],seed[2994],seed[63],seed[3359],seed[2043],seed[66],seed[534],seed[3217],seed[2012],seed[1208],seed[1313],seed[2432],seed[2297],seed[3197],seed[651],seed[729],seed[1870],seed[459],seed[374],seed[3491],seed[1468],seed[2339],seed[3011],seed[1754],seed[3533],seed[457],seed[2672],seed[1341],seed[781],seed[3354],seed[780],seed[2459],seed[1276],seed[3127],seed[3313],seed[632],seed[3766],seed[853],seed[206],seed[2762],seed[1873],seed[1655],seed[963],seed[2463],seed[2511],seed[718],seed[2033],seed[1865],seed[896],seed[4084],seed[851],seed[1549],seed[1302],seed[3094],seed[608],seed[2294],seed[1159],seed[3452],seed[2499],seed[3511],seed[1670],seed[3315],seed[1268],seed[342],seed[1255],seed[3535],seed[3121],seed[563],seed[997],seed[738],seed[2262],seed[1400],seed[1196],seed[3496],seed[200],seed[210],seed[3660],seed[3852],seed[2298],seed[2835],seed[1770],seed[1906],seed[2858],seed[419],seed[3264],seed[2588],seed[3270],seed[477],seed[2250],seed[1952],seed[3189],seed[3229],seed[1695],seed[1829],seed[3258],seed[3320],seed[452],seed[14],seed[978],seed[222],seed[2445],seed[3446],seed[918],seed[1516],seed[3685],seed[672],seed[3795],seed[2690],seed[3974],seed[2854],seed[3097],seed[188],seed[1652],seed[1024],seed[3584],seed[964],seed[285],seed[1650],seed[1984],seed[1712],seed[2747],seed[1121],seed[2875],seed[3478],seed[1942],seed[2242],seed[1493],seed[3782],seed[2389],seed[2521],seed[971],seed[2076],seed[488],seed[3269],seed[952],seed[3894],seed[2497],seed[1948],seed[2068],seed[2609],seed[3891],seed[3783],seed[3861],seed[3585],seed[3199],seed[2617],seed[2161],seed[2356],seed[1734],seed[2164],seed[4072],seed[253],seed[824],seed[2519],seed[600],seed[3445],seed[3272],seed[2042],seed[503],seed[3730],seed[443],seed[4085],seed[3343],seed[3404],seed[1735],seed[3221],seed[3798],seed[3560],seed[3658],seed[47],seed[903],seed[2373],seed[2999],seed[2611],seed[857],seed[3486],seed[1348],seed[3167],seed[3615],seed[3530],seed[2400],seed[1342],seed[558],seed[3365],seed[2248],seed[3529],seed[838],seed[3400],seed[435],seed[3880],seed[3295],seed[2132],seed[1358],seed[3960],seed[4022],seed[2985],seed[3757],seed[763],seed[2901],seed[1499],seed[2638],seed[2343],seed[2992],seed[1198],seed[3071],seed[65],seed[2119],seed[256],seed[2268],seed[646],seed[1308],seed[1144],seed[2558],seed[3661],seed[3752],seed[340],seed[931],seed[771],seed[2549],seed[106],seed[4054],seed[2413],seed[2310],seed[1298],seed[3555],seed[1262],seed[1737],seed[3634],seed[1047],seed[2289],seed[3517],seed[1114],seed[1854],seed[80],seed[634],seed[2867],seed[846],seed[3649],seed[766],seed[3561],seed[3854],seed[3025],seed[3012],seed[3727],seed[2073],seed[658],seed[3509],seed[3628],seed[2731],seed[3886],seed[2853],seed[2898],seed[299],seed[2648],seed[752],seed[1464],seed[3169],seed[3218],seed[1710],seed[1322],seed[29],seed[4042],seed[1123],seed[3970],seed[368],seed[3984],seed[2504],seed[756],seed[3226],seed[1885],seed[2473],seed[1469],seed[298],seed[2141],seed[2576],seed[3856],seed[553],seed[1133],seed[580],seed[1393],seed[3659],seed[3613],seed[3168],seed[2088],seed[4094],seed[3000],seed[1370],seed[1146],seed[751],seed[2290],seed[3402],seed[152],seed[26],seed[2426],seed[3729],seed[2282],seed[1796],seed[3116],seed[707],seed[2158],seed[1623],seed[1925],seed[3069],seed[3041],seed[3441],seed[2972],seed[2626],seed[3709],seed[3472],seed[1647],seed[1437],seed[2779],seed[1904],seed[3914],seed[906],seed[105],seed[333],seed[3952],seed[3991],seed[2360],seed[3859],seed[1544],seed[955],seed[736],seed[3497],seed[1245],seed[1264],seed[55],seed[1244],seed[576],seed[4089],seed[2085],seed[2701],seed[1964],seed[381],seed[427],seed[3677],seed[1908],seed[1278],seed[3583],seed[1092],seed[2124],seed[3484],seed[190],seed[2107],seed[2181],seed[2932],seed[863],seed[2730],seed[2514],seed[1174],seed[3463],seed[2218],seed[557],seed[1926],seed[4032],seed[3487],seed[885],seed[3872],seed[3995],seed[120],seed[2197],seed[3640],seed[2361],seed[231],seed[2450],seed[1768],seed[3345],seed[509],seed[2897],seed[4091],seed[620],seed[19],seed[297],seed[1501],seed[631],seed[996],seed[1922],seed[117],seed[2386],seed[1741],seed[2584],seed[3067],seed[1588],seed[2196],seed[1830],seed[2515],seed[2154],seed[1511],seed[2293],seed[3701],seed[3245],seed[3899],seed[900],seed[2996],seed[2675],seed[2964],seed[1211],seed[1147],seed[1087],seed[2163],seed[2175],seed[3163],seed[1913],seed[3302],seed[1131],seed[3896],seed[539],seed[679],seed[3776],seed[1386],seed[2900],seed[486],seed[2031],seed[1136],seed[2030],seed[2751],seed[3347],seed[216],seed[4050],seed[1299],seed[2995],seed[3637],seed[2337],seed[146],seed[2772],seed[103],seed[3526],seed[1574],seed[929],seed[3616],seed[3483],seed[3394],seed[2442],seed[1895],seed[2843],seed[827],seed[335],seed[3085],seed[2891],seed[148],seed[1746],seed[1852],seed[1832],seed[3372],seed[1941],seed[1072],seed[1484],seed[1070],seed[1568],seed[3066],seed[652],seed[1032],seed[841],seed[3608],seed[1801],seed[882],seed[1241],seed[1195],seed[1855],seed[1965],seed[3550],seed[3905],seed[2698],seed[362],seed[2699],seed[2317],seed[1170],seed[3287],seed[1557],seed[3206],seed[1728],seed[3519],seed[3430],seed[1532],seed[2465],seed[3309],seed[828],seed[3883],seed[3840],seed[1792],seed[487],seed[516],seed[165],seed[2899],seed[2967],seed[3948],seed[3170],seed[1073],seed[2629],seed[2251],seed[13],seed[2802],seed[2688],seed[607],seed[689],seed[1939],seed[949],seed[659],seed[3024],seed[1316],seed[1985],seed[999],seed[811],seed[4071],seed[2870],seed[350],seed[782],seed[423],seed[2712],seed[1398],seed[3062],seed[496],seed[1200],seed[69],seed[2436],seed[3393],seed[3339],seed[149],seed[965],seed[3209],seed[1215],seed[531],seed[3275],seed[3676],seed[1867],seed[586],seed[3621],seed[1857],seed[674],seed[2968],seed[1766],seed[2487],seed[3668],seed[945],seed[1573],seed[1366],seed[2502],seed[4045],seed[3707],seed[1793],seed[1292],seed[3458],seed[476],seed[3420],seed[2764],seed[1809],seed[2949],seed[988],seed[1296],seed[2903],seed[1321],seed[1183],seed[3188],seed[3379],seed[1699],seed[2257],seed[761],seed[193],seed[1752],seed[1896],seed[2274],seed[191],seed[3983],seed[3841],seed[283],seed[1848],seed[1745],seed[1052],seed[861],seed[2344],seed[3325],seed[732],seed[2071],seed[139],seed[1150],seed[3645],seed[3134],seed[425],seed[3811],seed[1633],seed[2002],seed[995],seed[2976],seed[795],seed[3579],seed[2546],seed[874],seed[182],seed[3407],seed[3712],seed[2615],seed[3527],seed[3408],seed[624],seed[3010],seed[2633],seed[623],seed[1161],seed[2346],seed[2890],seed[301],seed[1894],seed[1345],seed[426],seed[3459],seed[410],seed[2434],seed[1335],seed[3279],seed[1225],seed[2785],seed[643],seed[3961],seed[2823],seed[3946],seed[3182],seed[2482],seed[2377],seed[2309],seed[3962],seed[3166],seed[3026],seed[3557],seed[2709],seed[681],seed[1109],seed[1141],seed[2050],seed[726],seed[2708],seed[3719],seed[1337],seed[2622],seed[1617],seed[3630],seed[167],seed[1664],seed[33],seed[3351],seed[1062],seed[3745],seed[511],seed[3830],seed[3457],seed[2736],seed[1424],seed[1928],seed[1387],seed[324],seed[1786],seed[1272],seed[2117],seed[3323],seed[2249],seed[3534],seed[2906],seed[1003],seed[2078],seed[3439],seed[2077],seed[2643],seed[3870],seed[168],seed[3687],seed[237],seed[992],seed[4002],seed[1654],seed[1325],seed[589],seed[1307],seed[2475],seed[3185],seed[2391],seed[2657],seed[205],seed[2004],seed[3796],seed[3043],seed[3036],seed[1392],seed[1478],seed[1740],seed[556],seed[1524],seed[847],seed[3626],seed[2902],seed[1899],seed[2563],seed[3399],seed[404],seed[246],seed[3818],seed[3409],seed[3376],seed[1651],seed[3747],seed[71],seed[1555],seed[1911],seed[1760],seed[282],seed[719],seed[3921],seed[454],seed[1600],seed[3479],seed[341],seed[264],seed[258],seed[1982],seed[2203],seed[3032],seed[3001],seed[1045],seed[3710],seed[602],seed[2061],seed[2583],seed[2474],seed[3777],seed[3629],seed[2864],seed[533],seed[1636],seed[2811],seed[135],seed[2469],seed[926],seed[891],seed[1730],seed[2654],seed[378],seed[2569],seed[1005],seed[1056],seed[3361],seed[1021],seed[123],seed[275],seed[88],seed[2205],seed[3528],seed[1738],seed[2828],seed[3773],seed[987],seed[555],seed[639],seed[1759],seed[3797],seed[4065],seed[3341],seed[3505],seed[1627],seed[2941],seed[3332],seed[1637],seed[981],seed[2522],seed[2246],seed[609],seed[116],seed[1667],seed[1990],seed[3378],seed[2086],seed[1465],seed[3215],seed[1621],seed[1969],seed[2800],seed[2926],seed[1630],seed[2750],seed[2732],seed[2610],seed[3122],seed[377],seed[2278],seed[2340],seed[3271],seed[1490],seed[3058],seed[3577],seed[1135],seed[384],seed[2997],seed[3383],seed[2122],seed[3037],seed[1715],seed[3609],seed[3057],seed[3211],seed[2632],seed[1180],seed[3778],seed[1285],seed[2481],seed[1175],seed[3240],seed[4008],seed[85],seed[1860],seed[1962],seed[1641],seed[3410],seed[3698],seed[3280],seed[3002],seed[3562],seed[1644],seed[2943],seed[2462],seed[471],seed[585],seed[2556],seed[3614],seed[107],seed[2861],seed[1696],seed[1560],seed[2669],seed[2496],seed[352],seed[1596],seed[2880],seed[1584],seed[4043],seed[1129],seed[2857],seed[393],seed[3329],seed[1878],seed[597],seed[2051],seed[1126],seed[1886],seed[3088],seed[3089],seed[2108],seed[1826],seed[2946],seed[2005],seed[2774],seed[1811],seed[2001],seed[2939],seed[1638],seed[2191],seed[173],seed[1328],seed[875],seed[913],seed[2815],seed[749],seed[1933],seed[3131],seed[3101],seed[1818],seed[3785],seed[2984],seed[178],seed[1893],seed[1054],seed[1412],seed[445],seed[3741],seed[490],seed[3391],seed[3267],seed[217],seed[37],seed[3784],seed[1429],seed[2630],seed[4049],seed[1679],seed[230],seed[1601],seed[1267],seed[2238],seed[3780],seed[3909],seed[2171],seed[3114],seed[1452],seed[2507],seed[3596],seed[3824],seed[3823],seed[1678],seed[227],seed[28],seed[3652],seed[3423],seed[2613],seed[166],seed[2908],seed[1749],seed[2553],seed[3429],seed[572],seed[3130],seed[3033],seed[344],seed[1001],seed[1079],seed[1782],seed[3319],seed[3930],seed[1502],seed[3969],seed[2003],seed[2415],seed[2026],seed[1781],seed[627],seed[1026],seed[3646],seed[656],seed[3009],seed[1360],seed[3413],seed[541],seed[3926],seed[1645],seed[2069],seed[2328],seed[197],seed[2451],seed[3139],seed[2577],seed[3839],seed[2098],seed[1937],seed[2279],seed[1838],seed[1890],seed[938],seed[723],seed[3832],seed[787],seed[3427],seed[429],seed[4056],seed[912],seed[1237],seed[1098],seed[919],seed[954],seed[3181],seed[1841],seed[3187],seed[3506],seed[2850],seed[1763],seed[785],seed[3672],seed[3330],seed[2199],seed[1872],seed[2683],seed[2148],seed[794],seed[1102],seed[1534],seed[2215],seed[3688],seed[1018],seed[768],seed[1739],seed[3768],seed[1543],seed[300],seed[1000],seed[3897],seed[1779],seed[3428],seed[3165],seed[3695],seed[969],seed[2682],seed[3788],seed[3931],seed[4063],seed[986],seed[1954],seed[692],seed[3406],seed[3553],seed[3549],seed[1971],seed[1869],seed[917],seed[3792],seed[402],seed[1577],seed[1293],seed[2716],seed[367],seed[933],seed[665],seed[372],seed[1023],seed[2580],seed[3142],seed[1955],seed[4090],seed[343],seed[1152],seed[2485],seed[3495],seed[1720],seed[1592],seed[1140],seed[2168],seed[3989],seed[3806],seed[1431],seed[748],seed[2054],seed[1874],seed[1363],seed[2027],seed[543],seed[3851],seed[305],seed[3543],seed[83],seed[3597],seed[3091],seed[2425],seed[3665],seed[3431],seed[770],seed[1067],seed[2678],seed[1918],seed[3308],seed[2363],seed[1414],seed[4016],seed[3135],seed[104],seed[2844],seed[1265],seed[1691],seed[4014],seed[3070],seed[2492],seed[1483],seed[3935],seed[3760],seed[3019],seed[2767],seed[3641],seed[391],seed[2052],seed[3433],seed[3518],seed[3369],seed[1488],seed[357],seed[2631],seed[2149],seed[1665],seed[1317],seed[2285],seed[428],seed[3230],seed[3751],seed[760],seed[813],seed[3054],seed[240],seed[2303],seed[2754],seed[127],seed[112],seed[1344],seed[169],seed[1350],seed[549],seed[223],seed[271],seed[3395],seed[2595],seed[409],seed[3900],seed[2667],seed[2889],seed[662],seed[1275],seed[2572],seed[2190],seed[2133],seed[4093],seed[304],seed[613],seed[626],seed[1716],seed[3455],seed[3490],seed[1286],seed[2784],seed[517],seed[2973],seed[2495],seed[592],seed[3076],seed[2048],seed[2449],seed[1381],seed[3539],seed[848],seed[126],seed[3732],seed[2049],seed[1297],seed[1615],seed[3387],seed[1987],seed[1356],seed[705],seed[3653],seed[411],seed[1772],seed[61],seed[1230],seed[2437],seed[3034],seed[2381],seed[582],seed[1154],seed[128],seed[2816],seed[2269],seed[3064],seed[3655],seed[3086],seed[243],seed[2130],seed[336],seed[311],seed[618],seed[1042],seed[3889],seed[1940],seed[2228],seed[1821],seed[158],seed[2292],seed[1034],seed[1718],seed[3177],seed[2471],seed[856],seed[1055],seed[849],seed[2618],seed[2466],seed[2333],seed[279],seed[115],seed[973],seed[96],seed[3631],seed[1082],seed[3128],seed[880],seed[3467],seed[3397],seed[1213],seed[265],seed[3620],seed[1132],seed[650],seed[1086],seed[2147],seed[561],seed[2349],seed[291],seed[1572],seed[2684],seed[3713],seed[347],seed[2256],seed[1970],seed[1492],seed[3237],seed[817],seed[2813],seed[2888],seed[4035],seed[194],seed[2134],seed[327],seed[3462],seed[1866],seed[2272],seed[3642],seed[2179],seed[1404],seed[3243],seed[1256],seed[1812],seed[1188],seed[2725],seed[2390],seed[3794],seed[1435],seed[2804],seed[907],seed[184],seed[734],seed[1015],seed[3007],seed[2752],seed[3865],seed[1112],seed[3636],seed[3375],seed[2411],seed[461],seed[1145],seed[2165],seed[1642],seed[3567],seed[2029],seed[1331],seed[2245],seed[943],seed[4067],seed[3384],seed[1074],seed[2484],seed[3647],seed[108],seed[1871],seed[2616],seed[3589],seed[1512],seed[3895],seed[2221],seed[2925],seed[437],seed[3702],seed[2554],seed[2423],seed[3761],seed[1708],seed[3077],seed[4051],seed[2393],seed[737],seed[2448],seed[1729],seed[358],seed[1656],seed[379],seed[2776],seed[3986],seed[2345],seed[491],seed[1515],seed[2498],seed[953],seed[2532],seed[3083],seed[3913],seed[829],seed[524],seed[2733],seed[3749],seed[3575],seed[1542],seed[2186],seed[1011],seed[823],seed[1936],seed[2100],seed[3881],seed[2302],seed[1427],seed[1261],seed[453],seed[4001],seed[185],seed[960],seed[830],seed[1007],seed[741],seed[189],seed[415],seed[1269],seed[17],seed[254],seed[434],seed[1081],seed[1802],seed[1326],seed[442],seed[67],seed[2311],seed[2072],seed[1458],seed[2860],seed[1059],seed[1593],seed[2022],seed[833],seed[1446],seed[444],seed[2605],seed[1517],seed[212],seed[1038],seed[3079],seed[3153],seed[1153],seed[3968],seed[3787],seed[2674],seed[4],seed[1433],seed[288],seed[276],seed[3065],seed[1657],seed[1457],seed[909],seed[2797],seed[869],seed[406],seed[3082],seed[1439],seed[2483],seed[2905],seed[337],seed[225],seed[1823],seed[3039],seed[968],seed[816],seed[2472],seed[201],seed[1362],seed[3255],seed[1138],seed[2307],seed[696],seed[302],seed[1496],seed[717],seed[1778],seed[2722],seed[1530],seed[2713],seed[90],seed[3835],seed[686],seed[1916],seed[3965],seed[515],seed[2952],seed[1947],seed[868],seed[1085],seed[176],seed[3893],seed[3678],seed[3492],seed[750],seed[1595],seed[1807],seed[3820],seed[1380],seed[2944],seed[1221],seed[722],seed[4088],seed[53],seed[2718],seed[403],seed[560],seed[4044],seed[1078],seed[1019],seed[2461],seed[860],seed[1020],seed[3838],seed[892],seed[2136],seed[1388],seed[1727],seed[3277],seed[680],seed[2229],seed[2527],seed[500],seed[1039],seed[2545],seed[1960],seed[1538],seed[1634],seed[2167],seed[2503],seed[1181],seed[1725],seed[1139],seed[2661],seed[2145],seed[1688],seed[1201],seed[1546],seed[3117],seed[2934],seed[2429],seed[3759],seed[3016],seed[3172],seed[759],seed[3418],seed[685],seed[2300],seed[2094],seed[1923],seed[3074],seed[2839],seed[187],seed[859],seed[902],seed[805],seed[3417],seed[1455],seed[3919],seed[2446],seed[3541],seed[3502],seed[1049],seed[3202],seed[1723],seed[2101],seed[3132],seed[1119],seed[2988],seed[1474],seed[130],seed[2574],seed[2548],seed[2991],seed[611],seed[35],seed[972],seed[835],seed[3592],seed[2367],seed[48],seed[1158],seed[3224],seed[1162],seed[2066],seed[1258],seed[2827],seed[3936],seed[3618],seed[2110],seed[2517],seed[1755],seed[2539],seed[3885],seed[3364],seed[4046],seed[2371],seed[1002],seed[2477],seed[3873],seed[3573],seed[3042],seed[2277],seed[2612],seed[2280],seed[3736],seed[3092],seed[837],seed[4070],seed[2916],seed[2918],seed[3355],seed[2960],seed[366],seed[2129],seed[744],seed[3610],seed[2045],seed[588],seed[3363],seed[1312],seed[2213],seed[1339],seed[4020],seed[3254],seed[3027],seed[351],seed[1988],seed[2938],seed[1184],seed[3571],seed[2506],seed[1359],seed[2571],seed[1620],seed[2304],seed[2422],seed[363],seed[3450],seed[3476],seed[521],seed[2881],seed[2769],seed[776],seed[1856],seed[75],seed[767],seed[2935],seed[274],seed[1064],seed[1619],seed[2464],seed[1639],seed[125],seed[2872],seed[1476],seed[1974],seed[3971],seed[2760],seed[826],seed[289],seed[1846],seed[1762],seed[697],seed[803],seed[1669],seed[801],seed[345],seed[3808],seed[3774],seed[1677],seed[2805],seed[2338],seed[3356],seed[1521],seed[2636],seed[1949],seed[3102],seed[644],seed[2399],seed[1352],seed[323],seed[3120],seed[3673],seed[3699],seed[2385],seed[2624],seed[1487],seed[209],seed[1649],seed[3198],seed[3358],seed[1330],seed[2755],seed[4003],seed[598],seed[481],seed[2222],seed[1525],seed[3957],seed[2707],seed[1514],seed[4005],seed[1683],seed[2234],seed[2267],seed[731],seed[3157],seed[3105],seed[671],seed[3876],seed[1858],seed[181],seed[1658],seed[552],seed[3680],seed[2143],seed[3396],seed[655],seed[2808],seed[4057],seed[3008],seed[1430],seed[1950],seed[180],seed[786],seed[450],seed[2884],seed[260],seed[2728],seed[1413],seed[706],seed[2187],seed[2146],seed[499],seed[1409],seed[1438],seed[316],seed[1410],seed[3314],seed[2288],seed[1014],seed[1378],seed[3412],seed[1205],seed[1220],seed[204],seed[1450],seed[3328],seed[4095],seed[2478],seed[98],seed[1897],seed[2324],seed[473],seed[2153],seed[2336],seed[2568],seed[2526],seed[3906],seed[3246],seed[3178],seed[3624],seed[1537],seed[3866],seed[420],seed[3836],seed[1217],seed[4073],seed[1721],seed[3180],seed[538],seed[3235],seed[3371],seed[3090],seed[3878],seed[2118],seed[49],seed[3453],seed[1567],seed[2264],seed[3104],seed[1690],seed[2253],seed[495],seed[3635],seed[3879],seed[3548],seed[3063],seed[1029],seed[1847],seed[1605],seed[1709],seed[510],seed[2543],seed[742],seed[2642],seed[2489],seed[1840],seed[2299],seed[975],seed[2123],seed[2695],seed[3435],seed[603],seed[3800],seed[799],seed[698],seed[1461],seed[3093],seed[2687],seed[1612],seed[3939],seed[1684],seed[3059],seed[396],seed[4077],seed[1570],seed[2470],seed[3190],seed[383],seed[2192],seed[1017],seed[2057],seed[1836],seed[2789],seed[244],seed[3993],seed[2216],seed[3331],seed[2570],seed[174],seed[1790],seed[3964],seed[2676],seed[2510],seed[3918],seed[1240],seed[2034],seed[1518],seed[2693],seed[3547],seed[2178],seed[380],seed[2064],seed[3607],seed[898],seed[4087],seed[2301],seed[2263],seed[77],seed[962],seed[548],seed[1536],seed[2270],seed[1475],seed[431],seed[1309],seed[4011],seed[1310],seed[132],seed[1602],seed[2056],seed[529],seed[4017],seed[1130],seed[1685],seed[3718],seed[4026],seed[1613],seed[1459],seed[3988],seed[3151],seed[3942],seed[3256],seed[3985],seed[2023],seed[2070],seed[1610],seed[502],seed[1726],seed[4021],seed[1374],seed[3941],seed[467],seed[1440],seed[3155],seed[56],seed[2041],seed[3531],seed[3040],seed[940],seed[1243],seed[4025],seed[242],seed[1785],seed[3587],seed[1861],seed[2160],seed[2308],seed[2018],seed[3693],seed[1473],seed[1191],seed[3003],seed[873],seed[1384],seed[668],seed[91],seed[2724],seed[213],seed[136],seed[3179],seed[2537],seed[3588],seed[3306],seed[134],seed[3536],seed[4031],seed[3576],seed[4013],seed[4034],seed[2112],seed[3770],seed[2276],seed[1736],seed[1673],seed[2325],seed[2185],seed[334],seed[1389],seed[1853],seed[2865],seed[1168],seed[730],seed[1758],seed[930],seed[2347],seed[2096],seed[1445],seed[3436],seed[3061],seed[3119],seed[3029],seed[1761],seed[1824],seed[3191],seed[2099],seed[2882],seed[3554],seed[1010],seed[1422],seed[3847],seed[2673],seed[145],seed[1037],seed[814],seed[3447],seed[418],seed[2362],seed[1814],seed[1986],seed[2488],seed[2544],seed[2555],seed[3161],seed[695],seed[3803],seed[3513],seed[743],seed[57],seed[3096],seed[1122],seed[113],seed[879],seed[666],seed[1343],seed[3103],seed[3683],seed[2523],seed[400],seed[2706],seed[3756],seed[198],seed[1868],seed[594],seed[3299],seed[3485],seed[514],seed[3692],seed[1295],seed[1165],seed[571],seed[318],seed[2766],seed[716],seed[3723],seed[1113],seed[3944],seed[2711],seed[3437],seed[1753],seed[3917],seed[4030],seed[3377],seed[1320],seed[3304],seed[2501],seed[765],seed[1907],seed[464],seed[2468],seed[2159],seed[2162],seed[3972],seed[3663],seed[3137],seed[1234],seed[3604],seed[1912],seed[724],seed[1282],seed[4010],seed[1364],seed[806],seed[2180],seed[2177],seed[2691],seed[1794],seed[482],seed[3263],seed[43],seed[1609],seed[1110],seed[2271],seed[660],seed[2540],seed[164],seed[3149],seed[2876],seed[4038],seed[2749],seed[2443],seed[3186],seed[1917],seed[1226],seed[1303],seed[1382],seed[4083],seed[3247],seed[3725],seed[1978],seed[3799],seed[1663],seed[1963],seed[1661],seed[1173],seed[3389],seed[1084],seed[2379],seed[1548],seed[1581],seed[2140],seed[86],seed[2139],seed[1631],seed[1565],seed[1016],seed[3857],seed[1662],seed[669],seed[2593],seed[2235],seed[493],seed[1556],seed[3643],seed[1827],seed[203],seed[2971],seed[1882],seed[2573],seed[2729],seed[3388],seed[1008],seed[1820],seed[2105],seed[1604],seed[2286],seed[469],seed[2182],seed[1481],seed[1498],seed[3714],seed[1120],seed[2681],seed[821],seed[2457],seed[2369],seed[2830],seed[2841],seed[192],seed[3949],seed[2380],seed[3654],seed[2152],seed[788],seed[62],seed[424],seed[1945],seed[3537],seed[2174],seed[121],seed[1731],seed[1769],seed[2024],seed[4028],seed[779],seed[3500],seed[3095],seed[1338],seed[2792],seed[3568],seed[2220],seed[294],seed[3259],seed[3580],seed[2966],seed[3469],seed[2224],seed[593],seed[2259],seed[163],seed[4029],seed[89],seed[635],seed[2814],seed[1648],seed[3664],seed[1686],seed[501],seed[2028],seed[2644],seed[3367],seed[398],seed[179],seed[4036],seed[2114],seed[2700],seed[1681],seed[2211],seed[1124],seed[218],seed[961],seed[1603],seed[1576],seed[4033],seed[32],seed[1810],seed[710],seed[1523],seed[3081],seed[2538],seed[3769],seed[1036],seed[2254],seed[331],seed[619],seed[1747],seed[1231],seed[916],seed[2810],seed[670],seed[2856],seed[2909],seed[2989],seed[3833],seed[1552],seed[1875],seed[3657],seed[153],seed[1887],seed[2845],seed[2189],seed[2396],seed[119],seed[1247],seed[2258],seed[1239],seed[897],seed[1167],seed[27],seed[2352],seed[1732],seed[1668],seed[4079],seed[866],seed[376],seed[280],seed[3570],seed[224],seed[2109],seed[64],seed[2634],seed[764],seed[1733],seed[401],seed[3392],seed[2799],seed[2252],seed[3370],seed[1694],seed[663],seed[2102],seed[3650],seed[1171],seed[715],seed[2355],seed[4000],seed[1403],seed[1327],seed[2419],seed[1192],seed[3176],seed[3118],seed[4061],seed[667],seed[2956],seed[1594],seed[292],seed[3348],seed[2010],seed[2866],seed[2979],seed[2015],seed[3625],seed[3285],seed[3087],seed[2715],seed[3281],seed[546],seed[974],seed[1372],seed[438],seed[82],seed[3257],seed[1209],seed[1608],seed[1563],seed[3746],seed[758],seed[991],seed[40],seed[1539],seed[2798],seed[259],seed[1223],seed[2770],seed[3704],seed[3516],seed[1236],seed[2855],seed[2366],seed[3503],seed[3380],seed[2322],seed[1190],seed[78],seed[3262],seed[2414],seed[2565],seed[295],seed[2977],seed[2237],seed[527],seed[3786],seed[605],seed[2887],seed[1118],seed[3312],seed[1104],seed[2788],seed[1995],seed[3738],seed[3473],seed[494],seed[1803],seed[440],seed[1513],seed[746],seed[628],seed[177],seed[1428],seed[1509],seed[1194],seed[2201],seed[329],seed[2209],seed[574],seed[2067],seed[3470],seed[3563],seed[4068],seed[834],seed[3703],seed[775],seed[485],seed[1324],seed[322],seed[3239],seed[836],seed[3638],seed[30],seed[303],seed[45],seed[2852],seed[542],seed[944],seed[1629],seed[721],seed[2327],seed[2062],seed[1611],seed[2359],seed[1479],seed[3241],seed[862],seed[3812],seed[1956],seed[649],seed[793],seed[596],seed[2508],seed[1164],seed[3078],seed[2778],seed[899],seed[3159],seed[3674],seed[1186],seed[2312],seed[1800],seed[1780],seed[1806],seed[478],seed[1813],seed[142],seed[2692],seed[1898],seed[371],seed[3932],seed[2372],seed[3424],seed[1248],seed[2090],seed[31],seed[1957],seed[3223],seed[2316],seed[1116],seed[2833],seed[4059],seed[1616],seed[1289],seed[2331],seed[3073],seed[3816],seed[1701],seed[1526],seed[508],seed[1462],seed[2986],seed[3493],seed[2763],seed[2846],seed[3108],seed[3060],seed[364],seed[982],seed[2350],seed[3656],seed[2987],seed[3755],seed[1591],seed[1979],seed[2313],seed[1106],seed[2748],seed[1589],seed[599],seed[2421],seed[3566],seed[3871],seed[3353],seed[1408],seed[932],seed[3475],seed[2405],seed[3144],seed[3162],seed[439],seed[308],seed[2955],seed[3154],seed[2704],seed[23],seed[3877],seed[3922],seed[2019],seed[1825],seed[72],seed[1799],seed[1586],seed[1497],seed[893],seed[2040],seed[36],seed[16],seed[1053],seed[3236],seed[2886],seed[654],seed[519],seed[2155],seed[2607],seed[346],seed[818],seed[1334],seed[39],seed[831],seed[407],seed[1101],seed[1238],seed[309],seed[1697],seed[1281],seed[3868],seed[1561],seed[3422],seed[2226],seed[1724],seed[3310],seed[855],seed[622],seed[3763],seed[3194],seed[3822],seed[1176],seed[2740],seed[433],seed[3810],seed[2144],seed[518],seed[1227],seed[3052],seed[2374],seed[3411],seed[109],seed[1260],seed[284],seed[1347],seed[3220],seed[392],seed[3440],seed[1169],seed[1270],seed[1626],seed[1968],seed[645],seed[3244],seed[2579],seed[2032],seed[1336],seed[911],seed[2427],seed[1850],seed[3334],seed[2602],seed[1804],seed[1764],seed[2239],seed[979],seed[2975],seed[2650],seed[2600],seed[2877],seed[1961],seed[2231],seed[2831],seed[2121],seed[1012],seed[41],seed[233],seed[2341],seed[3338],seed[3288],seed[1551],seed[1880],seed[3775],seed[2589],seed[1743],seed[3669],seed[1383],seed[1905],seed[3827],seed[537],seed[2036],seed[3442],seed[310],seed[2458],seed[281],seed[2658],seed[1700],seed[3023],seed[3887],seed[884],seed[3099],seed[3115],seed[3234],seed[361],seed[399],seed[3013],seed[3265],seed[1319],seed[2726],seed[3726],seed[2416],seed[1357],seed[1066],seed[2980],seed[208],seed[1580],seed[3771],seed[3975],seed[52],seed[154],seed[3342],seed[2305],seed[3564],seed[2007],seed[1935],seed[547],seed[3924],seed[2335],seed[769],seed[1096],seed[3992],seed[1391],seed[920],seed[2320],seed[2969],seed[1043],seed[1099],seed[2490],seed[2874],seed[2170],seed[2598],seed[3521],seed[3021],seed[1271],seed[3336],seed[4053],seed[1989],seed[3860],seed[2],seed[590],seed[3599],seed[2561],seed[1822],seed[2758],seed[2065],seed[1547],seed[3603],seed[252],seed[3789],seed[1444],seed[1107],seed[1291],seed[1442],seed[2329],seed[456],seed[2398],seed[2401],seed[3344],seed[2623],seed[540],seed[2652],seed[3136],seed[1143],seed[3911],seed[1953],seed[3546],seed[1405],seed[38],seed[3686],seed[3595],seed[3350],seed[1103],seed[2008],seed[1578],seed[1419],seed[20],seed[3920],seed[2656],seed[3100],seed[1177],seed[2664],seed[3814],seed[3904],seed[155],seed[3742],seed[1235],seed[4069],seed[170],seed[2851],seed[3421],seed[390],seed[2097],seed[3477],seed[1900],seed[2686],seed[3508],seed[1006],seed[3123],seed[4023],seed[2592],seed[772],seed[3152],seed[3291],seed[277],seed[3862],seed[3826],seed[235],seed[3056],seed[1432],seed[263],seed[852],seed[3232],seed[871],seed[239],seed[3148],seed[1997],seed[2038],seed[262],seed[2358],seed[790],seed[1531],seed[832],seed[967],seed[161],seed[93],seed[858],seed[111],seed[840],seed[475],seed[985],seed[2645],seed[1973],seed[2225],seed[3700],seed[3606],seed[2440],seed[144],seed[2265],seed[3600],seed[3107],seed[3733],seed[3720],seed[3907],seed[3360],seed[3098],seed[483],seed[1454],seed[2564],seed[881],seed[4052],seed[621],seed[506],seed[800],seed[2476],seed[3804],seed[3160],seed[921],seed[1204],seed[889],seed[1575],seed[1083],seed[910],seed[2871],seed[3979],seed[701],seed[2993],seed[1750],seed[2382],seed[2207],seed[1839],seed[221],seed[1172],seed[3569],seed[1155],seed[42],seed[2803],seed[498],seed[1632],seed[3721],seed[1902],seed[3460],seed[50],seed[2275],seed[2486],seed[2849],seed[386],seed[397],seed[338],seed[2878],seed[2368],seed[234],seed[2394],seed[1467],seed[1914],seed[822],seed[2637],seed[54],seed[195],seed[1095],seed[5],seed[1706],seed[1022],seed[2697],seed[3126],seed[3416],seed[3201],seed[2281],seed[1128],seed[4041],seed[2868],seed[3138],seed[12],seed[1828],seed[1407],seed[2937],seed[1994],seed[983],seed[528],seed[2266],seed[2694],seed[1675],seed[3954],seed[1719],seed[2586],seed[2869],seed[2083],seed[1390],seed[1693],seed[3623],seed[2387],seed[2822],seed[2791],seed[3925],seed[3559],seed[3233],seed[2111],seed[630],seed[2365],seed[581],seed[1480],seed[3929],seed[1550],seed[1981],seed[1582],seed[3200],seed[2893],seed[739],seed[3212],seed[3357],seed[1643],seed[3910],seed[3133],seed[1314],seed[3207],seed[895],seed[2604],seed[2647],seed[3520],seed[3523],seed[1417],seed[2982],seed[802],seed[850],seed[1845],seed[3943],seed[2924],seed[2053],seed[2479],seed[2773],seed[939],seed[3959],seed[3020],seed[3203],seed[3278],seed[532],seed[2743],seed[2296],seed[653],seed[3110],seed[1704],seed[2370],seed[349],seed[2236],seed[266],seed[1698],seed[567],seed[2742],seed[3737],seed[3611],seed[3633],seed[2525],seed[507],seed[3174],seed[3675],seed[129],seed[3292],seed[990],seed[2444],seed[1274],seed[2092],seed[2198],seed[317],seed[914],seed[3927],seed[3289],seed[1938],seed[2156],seed[2208],seed[3648],seed[2663],seed[118],seed[4060],seed[1932],seed[2927],seed[942],seed[1773],seed[3318],seed[887],seed[1528],seed[545],seed[2826],seed[196],seed[3129],seed[1212],seed[2705],seed[2137],seed[1061],seed[2885],seed[2353],seed[2172],seed[1218],seed[791],seed[1862],seed[1711],seed[207],seed[3498],seed[3075],seed[4076],seed[1566],seed[3937],seed[784],seed[1351],seed[2079],seed[1713],seed[1206],seed[3875],seed[412],seed[3373],seed[2255],seed[2653],seed[3219],seed[1888],seed[577],seed[3684],seed[1368],seed[2035],seed[4082],seed[2084],seed[1406],seed[3143],seed[3048],seed[3915],seed[3482],seed[3958],seed[4075],seed[2786],seed[3158],seed[2670],seed[3779],seed[1756],seed[232],seed[601],seed[3337],seed[1263],seed[2765],seed[924],seed[1353],seed[711],seed[3728],seed[2157],seed[34],seed[2323],seed[44],seed[568],seed[3572],seed[2923],seed[51],seed[2491],seed[1471],seed[2717],seed[447],seed[708],seed[2668],seed[1046],seed[2200],seed[820],seed[1105],seed[1376],seed[2059],seed[3466],seed[1504],seed[2601],seed[2044],seed[3586],seed[1919],seed[808],seed[3109],seed[2796],seed[3928],seed[3767],seed[4080],seed[2737],seed[100],seed[2671],seed[1415],seed[2408],seed[3311],seed[1094],seed[1305],seed[2230],seed[1505],seed[2435],seed[465],seed[3781],seed[4009],seed[4086],seed[778],seed[2418],seed[640],seed[2500],seed[2025],seed[257],seed[2662],seed[2720],seed[267],seed[2582],seed[625],seed[2958],seed[3055],seed[2166],seed[3912],seed[1033],seed[3049],seed[2847],seed[3501],seed[1714],seed[3349],seed[1771],seed[3828],seed[1076],seed[3333],seed[3268],seed[584],seed[1004],seed[468],seed[1111],seed[2646],seed[1625],seed[2591],seed[682],seed[2424],seed[1117],seed[1495],seed[497],seed[890],seed[993],seed[2547],seed[610],seed[526],seed[472],seed[328],seed[865],seed[3544],seed[11],seed[3214],seed[2354],seed[3825],seed[87],seed[1795],seed[3031],seed[432],seed[2782],seed[1035],seed[1379],seed[1257],seed[21],seed[3558],seed[2665],seed[3346],seed[647],seed[1203],seed[946],seed[3015],seed[1125],seed[2516],seed[3791],seed[1411],seed[2227],seed[2006],seed[2921],seed[1399],seed[984],seed[3017],seed[3978],seed[3301],seed[2639],seed[3208],seed[220],seed[935],seed[3705],seed[1311],seed[3639],seed[3869],seed[2640],seed[566],seed[1687],seed[755],seed[365],seed[1569],seed[1722],seed[2840],seed[2961],seed[740],seed[559],seed[1214],seed[3374],seed[2914],seed[3303],seed[579],seed[796],seed[4004],seed[2524],seed[3973],seed[353],seed[479],seed[1876],seed[3340],seed[1646],seed[3205],seed[2428],seed[1808],seed[413],seed[612],seed[1443],seed[1606],seed[1744],seed[573],seed[3282],seed[2480],seed[2781],seed[1717],seed[1396],seed[3524],seed[332],seed[101],seed[3735],seed[713],seed[2575],seed[1983],seed[1819],seed[1929],seed[3963],seed[2628],seed[664],seed[2103],seed[725],seed[313],seed[1222],seed[2896],seed[3512],seed[1063],seed[3326],seed[2195],seed[2735],seed[1229],seed[2318],seed[2535],seed[4019],seed[421],seed[3171],seed[587],seed[2232],seed[4040],seed[249],seed[2635],seed[58],seed[3903],seed[2970],seed[306],seed[2357],seed[3853],seed[1931],seed[2453],seed[2193],seed[405],seed[1924],seed[3831],seed[637],seed[2873],seed[3204],seed[2513],seed[1520],seed[2000],seed[1494],seed[2509],seed[219],seed[2505],seed[3731],seed[1491],seed[3696],seed[1921],seed[94],seed[3790],seed[359],seed[4064],seed[356],seed[2917],seed[448],seed[1967],seed[2619],seed[2315],seed[2819],seed[1805],seed[449],seed[1508],seed[908],seed[3764],seed[1097],seed[1300],seed[512],seed[958],seed[1934],seed[360],seed[2689],seed[2913],seed[4074],seed[810],seed[2441],seed[1482],seed[1834],seed[774],seed[2406],seed[73],seed[894],seed[1323],seed[2074],seed[1423],seed[2801],seed[4039],seed[804],seed[97],seed[417],seed[575],seed[1776],seed[2562],seed[3793],seed[2397],seed[1607],seed[3252],seed[1426],seed[2095],seed[2859],seed[2702],seed[3849],seed[59],seed[2214],seed[3238],seed[1889],seed[3381],seed[617],seed[228],seed[1048],seed[904],seed[1702],seed[2392],seed[2787],seed[2395],seed[7],seed[2284],seed[3981],seed[1065],seed[1202],seed[261],seed[1242],seed[2212],seed[1028],seed[3140],seed[1506],seed[15],seed[131],seed[2587],seed[3716],seed[3815],seed[1210],seed[287],seed[520],seed[1127],seed[395],seed[2596],seed[1980],seed[684],seed[2243],seed[1185],seed[704],seed[2233],seed[2930],seed[2655],seed[1510],seed[1250],seed[3276],seed[1703],seed[1093],seed[1340],seed[3113],seed[1425],seed[905],seed[251],seed[2013],seed[797],seed[4062],seed[675],seed[3708],seed[3717],seed[1418],seed[2660],seed[2529],seed[3998],seed[1843],seed[3022],seed[1883],seed[3286],seed[3451],seed[4015],seed[3578],seed[2364],seed[2273],seed[2947],seed[3834],seed[1148],seed[2627],seed[3551],seed[3821],seed[1707],seed[3990],seed[642],seed[1901],seed[137],seed[46],seed[1585],seed[1],seed[138],seed[1972],seed[2106],seed[2247],seed[1705],seed[1587],seed[3322],seed[1903],seed[2039],seed[687],seed[451],seed[2135],seed[1628],seed[2848],seed[3867],seed[1998],seed[3327],seed[2542],seed[2082],seed[3722],seed[2978],seed[2614],seed[2824],seed[236],seed[1346],seed[484],seed[1108],seed[934],seed[1507],seed[877],seed[3997],seed[2780],seed[1013],seed[1775],seed[3405],seed[583],seed[2557],seed[2223],seed[901],seed[3807],seed[2113],seed[2836],seed[3976],seed[1365],seed[3266],seed[947],seed[3053],seed[922],seed[4037],seed[3293],seed[1249],seed[0],seed[2821],seed[354],seed[1069],seed[70],seed[3908],seed[2922],seed[1071],seed[76],seed[1777],seed[2863],seed[2757],seed[1672],seed[3898],seed[773],seed[2014],seed[888],seed[3951],seed[2680],seed[480],seed[1562],seed[2775],seed[2620],seed[3690],seed[1306],seed[2433],seed[3715],seed[1301],seed[3251],seed[677],seed[3739],seed[691],seed[2825],seed[319],seed[3662],seed[1666],seed[1598],seed[3581],seed[245],seed[2744],seed[2963],seed[314],seed[727],seed[387],seed[3845],seed[3858],seed[124],seed[4048],seed[3316],seed[4092],seed[114],seed[1394],seed[1676],seed[948],seed[604],seed[2104],seed[678],seed[1219],seed[68],seed[2910],seed[436],seed[2404],seed[3514],seed[3574],seed[1044],seed[1355],seed[2533],seed[1635],seed[1765],seed[2651],seed[3216],seed[3481],seed[133],seed[2291],seed[3454],seed[925],seed[339],seed[2009],seed[3748],seed[3438],seed[3863],seed[3283],seed[3605],seed[3744],seed[4066],seed[2016],seed[2528],seed[1590],seed[2998],seed[430],seed[733],seed[1246],seed[2438],seed[466],seed[286],seed[950],seed[513],seed[3632],seed[544],seed[3953],seed[2240],seed[2768],seed[1068],seed[2837],seed[1788],seed[3582],seed[1533],seed[2738],seed[3819],seed[1554],seed[2552],seed[700],seed[3471],seed[2384],seed[2531],seed[156],seed[3947],seed[2512],seed[422],seed[3260],seed[1266],seed[1944],seed[1653],seed[3499],seed[3601],seed[3444],seed[2021],seed[272],seed[3977],seed[4024],seed[2806],seed[1361],seed[4047],seed[2594],seed[3321],seed[3014],seed[2566],seed[1280],seed[2439],seed[3284],seed[2116],seed[3938],seed[3967],seed[1472],seed[569],seed[1091],seed[3125],seed[250],seed[3489],seed[325],seed[2940],seed[1774],seed[633],seed[815],seed[657],seed[1080],seed[3565],seed[1252],seed[3874],seed[2649],seed[2879],seed[2378],seed[1996],seed[2809],seed[1784],seed[2376],seed[385],seed[745],seed[1659],seed[3542],seed[2942],seed[388],seed[2334],seed[1863],seed[2075],seed[3305],seed[199],seed[3956],seed[3324],seed[3426],seed[1618],seed[636],seed[2741],seed[3192],seed[2794],seed[2807],seed[3261],seed[211],seed[3449],seed[2590],seed[226],seed[2974],seed[4027],seed[1436],seed[688],seed[1187],seed[2093],seed[886],seed[2017],seed[638],seed[1160],seed[1448],seed[3480],seed[3842],seed[2759],seed[3617],seed[505],seed[3227],seed[980],seed[3724],seed[1920],seed[183],seed[2559],seed[1891],seed[414],seed[3045],seed[1197],seed[215],seed[523],seed[3987],seed[1864],seed[702],seed[2115],seed[3671],seed[3890],seed[1682],seed[3864],seed[854],seed[3758],seed[3999],seed[348],seed[1660],seed[2260],seed[3667],seed[3106],seed[641],seed[1182],seed[9],seed[1851],seed[3390],seed[3196],seed[994],seed[1742],seed[2659],seed[151],seed[446],seed[1163],seed[3250],seed[3850],seed[845],seed[1149],seed[99],seed[3494],seed[535],seed[4055],seed[1142],seed[876],seed[2904],seed[2581],seed[2756],seed[728],seed[3141],seed[1692],seed[143],seed[1283],seed[798],seed[1030],seed[825],seed[1958],seed[3994],seed[2420],seed[10],seed[2011],seed[3150],seed[3050],seed[1304],seed[3934],seed[941],seed[186],seed[463],seed[1050],seed[1134],seed[3294],seed[870],seed[394],seed[3047],seed[1881],seed[3697],seed[3772],seed[24],seed[3461],seed[3147],seed[578],seed[735],seed[3743],seed[268],seed[1179],seed[753],seed[2409],seed[1842],seed[2818],seed[2920],seed[1915],seed[3044],seed[951],seed[2599],seed[2550],seed[1077],seed[2746],seed[3950],seed[3464],seed[2188],seed[3298],seed[3005],seed[355],seed[2244],seed[320],seed[2125],seed[3507],seed[3622],seed[2603],seed[1529],seed[290],seed[1031],seed[389],seed[1751],seed[2745],seed[3386],seed[3274],seed[1089],seed[1966],seed[616],seed[1354],seed[1976],seed[492],seed[1253],seed[1489],seed[160],seed[1318],seed[792],seed[1927],seed[2326],seed[2929],seed[147],seed[1477],seed[162],seed[2954],seed[2173],seed[2375],seed[1385],seed[757],seed[923],seed[3018],seed[699],seed[1100],seed[382],seed[3627],seed[3],seed[141],seed[3980],seed[2431],seed[293],seed[248],seed[1540],seed[3366],seed[3996],seed[1783],seed[2460],seed[3335],seed[883],seed[843],seed[1441],seed[842],seed[25],seed[3414],seed[3844],seed[1375],seed[4006],seed[2817],seed[977],seed[867],seed[122],seed[1402],seed[2951],seed[1456],seed[1470],seed[1519],seed[3515],seed[2892],seed[79],seed[3183],seed[1287],seed[1421],seed[1787],seed[3762],seed[2793],seed[3146],seed[1137],seed[3813],seed[2721],seed[3691],seed[525],seed[789],seed[1535],seed[998],seed[1193],seed[1930],seed[2518],seed[247],seed[1367],seed[844],seed[1156],seed[1259],seed[1434],seed[2907],seed[214],seed[2795],seed[1207],seed[3290],seed[1486],seed[1189],seed[375],seed[2089],seed[1377],seed[819],seed[2131],seed[2567],seed[315],seed[3228],seed[3945],seed[3030],seed[3368],seed[1559],seed[3072],seed[3802],seed[970],seed[3213],seed[2727],seed[2150],seed[1151],seed[2217],seed[2761],seed[2306],seed[3619],seed[3525],seed[812],seed[2965],seed[3809],seed[754],seed[709],seed[1789],seed[2194],seed[3432],seed[2151],seed[4018],seed[2953],seed[270],seed[458],seed[1397],seed[1251],seed[3694],seed[3175],seed[1288],seed[2219],seed[3242],seed[1597],seed[2883],seed[1835],seed[3902],seed[1041],seed[159],seed[1564],seed[1951],seed[460],seed[2832],seed[229],seed[1993],seed[3651],seed[3474],seed[81],seed[3124],seed[2931],seed[3385],seed[202],seed[3193],seed[2530],seed[330],seed[3173],seed[3038],seed[777],seed[959],seed[2060],seed[3545],seed[3916],seed[3888],seed[2447],seed[2342],seed[2402],seed[694],seed[2919],seed[1943],seed[1115],seed[2383],seed[1290],seed[1797],seed[3006],seed[3666],seed[2410],seed[321],seed[8],seed[4078],seed[1284],seed[3468],seed[2091],seed[3296],seed[1315],seed[1849],seed[1329],seed[2585],seed[1199],seed[3532],seed[2597],seed[2895],seed[2783],seed[1837],seed[976],seed[2981],seed[693],seed[84],seed[1815],seed[1216],seed[2241],seed[3594],seed[966],seed[2685],seed[1757],seed[3084],seed[554],seed[3843],seed[661],seed[370],seed[1332],seed[4012],seed[307],seed[1232],seed[3805],seed[2330],seed[3398],seed[3538],seed[489],seed[2834],seed[591],seed[1420],seed[1522],seed[3923],seed[570],seed[3248],seed[551],seed[470],seed[2541],seed[416],seed[2912],seed[1844],seed[3448],seed[2677],seed[326],seed[3164],seed[1485],seed[2842],seed[1859],seed[2838],seed[102],seed[3307],seed[3540],seed[937],seed[3754],seed[3382],seed[2606],seed[2204],seed[720],seed[1946],seed[4007],seed[2087],seed[2210],seed[2771],seed[3837],seed[1671],seed[783],seed[1090],seed[408],seed[3612],seed[2388],seed[3425],seed[2933],seed[1879],seed[3051],seed[2202],seed[2894],seed[2169],seed[2454],seed[3901],seed[3679],seed[2915],seed[690],seed[3882],seed[1553],seed[3955],seed[3552],seed[74],seed[3273],seed[1058],seed[1447],seed[172],seed[1401],seed[2412],seed[1009],seed[809],seed[3510],seed[2455],seed[3046],seed[3982],seed[3750],seed[3231],seed[2456],seed[2959],seed[872],seed[3415],seed[140],seed[1294],seed[1892],seed[2287],seed[175],seed[3035],seed[1909],seed[3184],seed[3644],seed[1224],seed[3401],seed[296],seed[369],seed[762],seed[683],seed[312],seed[1541],seed[3593],seed[3443],seed[3689],seed[1992],seed[1060],seed[564],seed[3456],seed[1624],seed[536],seed[3590],seed[1877],seed[278],seed[3765],seed[3682],seed[1831],seed[2957],seed[2348],seed[2493],seed[3711],seed[1166],seed[2127],seed[3300],seed[1767],seed[1527]}; 
//        seed9 <= {seed[260],seed[737],seed[3850],seed[3852],seed[2184],seed[422],seed[1938],seed[626],seed[753],seed[3877],seed[522],seed[4011],seed[60],seed[3657],seed[1669],seed[2945],seed[549],seed[1798],seed[3738],seed[2443],seed[2663],seed[2384],seed[851],seed[2015],seed[1088],seed[2265],seed[472],seed[1429],seed[1388],seed[2101],seed[3797],seed[3687],seed[946],seed[1090],seed[3151],seed[749],seed[262],seed[464],seed[747],seed[294],seed[3960],seed[672],seed[2219],seed[3893],seed[1908],seed[3924],seed[3750],seed[1568],seed[67],seed[3965],seed[3925],seed[1361],seed[536],seed[4084],seed[3574],seed[2701],seed[17],seed[820],seed[3895],seed[78],seed[2657],seed[2516],seed[321],seed[2159],seed[284],seed[392],seed[568],seed[2831],seed[1614],seed[2951],seed[1706],seed[3890],seed[1073],seed[1877],seed[1322],seed[771],seed[1256],seed[3918],seed[1271],seed[3961],seed[1081],seed[3222],seed[3365],seed[1895],seed[2475],seed[1520],seed[1664],seed[3744],seed[3701],seed[3772],seed[2827],seed[145],seed[1534],seed[223],seed[920],seed[3449],seed[4043],seed[1215],seed[2463],seed[3028],seed[2422],seed[230],seed[2494],seed[10],seed[1760],seed[2865],seed[2111],seed[1393],seed[1161],seed[3620],seed[3366],seed[871],seed[2260],seed[1855],seed[2414],seed[19],seed[4069],seed[3352],seed[1213],seed[1439],seed[1503],seed[163],seed[1363],seed[3896],seed[3052],seed[2278],seed[693],seed[1681],seed[526],seed[1595],seed[240],seed[809],seed[2526],seed[383],seed[2741],seed[1484],seed[2661],seed[2224],seed[80],seed[151],seed[1633],seed[2832],seed[1644],seed[1368],seed[832],seed[1165],seed[3327],seed[277],seed[3729],seed[1238],seed[416],seed[181],seed[1015],seed[2479],seed[106],seed[573],seed[3667],seed[810],seed[1834],seed[252],seed[1533],seed[2651],seed[3886],seed[484],seed[2131],seed[2783],seed[3487],seed[927],seed[1913],seed[1299],seed[2193],seed[382],seed[577],seed[118],seed[160],seed[1536],seed[2570],seed[2162],seed[479],seed[2069],seed[2989],seed[990],seed[1601],seed[3663],seed[1784],seed[2816],seed[2204],seed[3868],seed[2615],seed[885],seed[33],seed[2133],seed[2825],seed[3074],seed[1233],seed[1797],seed[1637],seed[4028],seed[2],seed[1435],seed[2129],seed[2499],seed[1096],seed[1738],seed[4068],seed[2503],seed[2396],seed[1675],seed[3742],seed[2483],seed[2359],seed[1773],seed[958],seed[3548],seed[1485],seed[1505],seed[1867],seed[3575],seed[2685],seed[1692],seed[3088],seed[9],seed[1655],seed[3811],seed[3810],seed[410],seed[2586],seed[1795],seed[3677],seed[2058],seed[1274],seed[760],seed[2904],seed[3529],seed[1513],seed[3482],seed[1626],seed[3038],seed[4080],seed[451],seed[698],seed[1310],seed[2502],seed[3165],seed[3872],seed[2141],seed[1323],seed[1390],seed[4021],seed[3361],seed[485],seed[2279],seed[2137],seed[3375],seed[1830],seed[2621],seed[3532],seed[1980],seed[3188],seed[1995],seed[714],seed[2839],seed[1351],seed[2815],seed[1979],seed[3398],seed[3658],seed[650],seed[2342],seed[2769],seed[489],seed[649],seed[2188],seed[1755],seed[1904],seed[121],seed[3261],seed[278],seed[3536],seed[1244],seed[783],seed[2729],seed[3702],seed[2256],seed[1703],seed[1756],seed[3335],seed[4083],seed[2763],seed[2361],seed[584],seed[2940],seed[1540],seed[1531],seed[2715],seed[811],seed[4085],seed[1075],seed[114],seed[1879],seed[854],seed[470],seed[3178],seed[2071],seed[1967],seed[2233],seed[4042],seed[1432],seed[2863],seed[3565],seed[1635],seed[2976],seed[476],seed[1964],seed[3061],seed[3369],seed[2728],seed[3220],seed[1340],seed[3092],seed[458],seed[2937],seed[2164],seed[667],seed[1001],seed[2477],seed[2762],seed[3413],seed[1929],seed[2196],seed[3539],seed[1229],seed[241],seed[1246],seed[1091],seed[957],seed[2946],seed[2488],seed[1876],seed[3740],seed[558],seed[2998],seed[1652],seed[1744],seed[882],seed[2645],seed[1304],seed[3727],seed[963],seed[3237],seed[1791],seed[92],seed[828],seed[2883],seed[3623],seed[887],seed[168],seed[499],seed[2474],seed[3119],seed[784],seed[2625],seed[1032],seed[2294],seed[4001],seed[3819],seed[3731],seed[726],seed[895],seed[245],seed[3224],seed[2211],seed[1611],seed[1321],seed[3],seed[388],seed[3194],seed[888],seed[3116],seed[3477],seed[1324],seed[3820],seed[3919],seed[994],seed[1739],seed[561],seed[1440],seed[542],seed[3948],seed[447],seed[2126],seed[3517],seed[1976],seed[1653],seed[563],seed[1122],seed[2482],seed[3084],seed[2374],seed[3436],seed[2817],seed[1730],seed[2529],seed[3757],seed[775],seed[3673],seed[1114],seed[2630],seed[567],seed[1647],seed[3916],seed[578],seed[3018],seed[2023],seed[425],seed[3577],seed[2844],seed[983],seed[1905],seed[2811],seed[3030],seed[759],seed[135],seed[1222],seed[4076],seed[3378],seed[3244],seed[1826],seed[2280],seed[2272],seed[3370],seed[3755],seed[681],seed[3037],seed[1582],seed[4022],seed[1207],seed[1950],seed[1766],seed[265],seed[3021],seed[1326],seed[655],seed[1139],seed[1620],seed[3474],seed[3480],seed[1731],seed[81],seed[2067],seed[2173],seed[2986],seed[2717],seed[2978],seed[3356],seed[2424],seed[1214],seed[4059],seed[3869],seed[2183],seed[2814],seed[2033],seed[2400],seed[841],seed[3763],seed[593],seed[3121],seed[270],seed[376],seed[3478],seed[2758],seed[1954],seed[924],seed[2476],seed[1859],seed[632],seed[24],seed[1226],seed[2754],seed[3271],seed[778],seed[3345],seed[1060],seed[3063],seed[3388],seed[870],seed[1374],seed[2478],seed[481],seed[1005],seed[2045],seed[3215],seed[452],seed[580],seed[620],seed[1162],seed[1003],seed[1259],seed[1893],seed[3911],seed[3341],seed[1850],seed[3706],seed[1423],seed[1287],seed[1919],seed[2667],seed[1884],seed[487],seed[3156],seed[740],seed[3445],seed[950],seed[3697],seed[1133],seed[2764],seed[1537],seed[1377],seed[2251],seed[2590],seed[930],seed[224],seed[3883],seed[1442],seed[1510],seed[674],seed[2709],seed[131],seed[1421],seed[2795],seed[562],seed[116],seed[507],seed[1254],seed[1932],seed[3363],seed[2725],seed[3389],seed[271],seed[2209],seed[285],seed[2680],seed[3636],seed[3174],seed[915],seed[772],seed[2852],seed[3837],seed[1205],seed[2270],seed[1914],seed[3198],seed[2934],seed[3241],seed[1977],seed[2489],seed[2267],seed[1722],seed[2583],seed[2650],seed[3679],seed[2303],seed[409],seed[3009],seed[3938],seed[3983],seed[2792],seed[492],seed[1149],seed[3200],seed[880],seed[897],seed[3932],seed[2580],seed[192],seed[362],seed[3034],seed[3199],seed[685],seed[3320],seed[724],seed[516],seed[1169],seed[607],seed[1425],seed[3471],seed[2659],seed[528],seed[2592],seed[4017],seed[1529],seed[3635],seed[3434],seed[1935],seed[1610],seed[3279],seed[3692],seed[389],seed[1911],seed[2755],seed[3977],seed[2149],seed[359],seed[253],seed[2076],seed[1196],seed[1695],seed[3336],seed[3264],seed[2561],seed[1105],seed[365],seed[3381],seed[4003],seed[341],seed[2991],seed[2740],seed[2223],seed[2089],seed[4053],seed[633],seed[328],seed[4044],seed[1415],seed[1183],seed[4012],seed[3722],seed[2871],seed[3280],seed[1565],seed[3934],seed[4052],seed[1912],seed[3286],seed[1454],seed[872],seed[1067],seed[2027],seed[2331],seed[611],seed[1062],seed[1087],seed[2026],seed[2834],seed[2555],seed[3664],seed[3616],seed[1378],seed[2077],seed[4073],seed[1843],seed[1632],seed[3380],seed[2882],seed[3265],seed[22],seed[1118],seed[1084],seed[764],seed[3631],seed[1143],seed[1469],seed[3659],seed[483],seed[2299],seed[1098],seed[1940],seed[3991],seed[2176],seed[1380],seed[2711],seed[3825],seed[105],seed[53],seed[838],seed[1209],seed[2011],seed[1342],seed[2138],seed[3922],seed[701],seed[1902],seed[1822],seed[2386],seed[1519],seed[3282],seed[3826],seed[3069],seed[3491],seed[2912],seed[1412],seed[3989],seed[503],seed[4078],seed[2720],seed[2132],seed[1587],seed[2339],seed[1414],seed[1251],seed[4082],seed[74],seed[3622],seed[3344],seed[873],seed[3598],seed[2369],seed[2050],seed[1449],seed[2212],seed[2931],seed[1642],seed[361],seed[457],seed[559],seed[2652],seed[1951],seed[3836],seed[3728],seed[1553],seed[3384],seed[218],seed[2771],seed[2363],seed[3470],seed[934],seed[411],seed[1943],seed[66],seed[85],seed[3259],seed[214],seed[101],seed[937],seed[1694],seed[3155],seed[3683],seed[2908],seed[1017],seed[3439],seed[3466],seed[4095],seed[736],seed[68],seed[490],seed[2139],seed[817],seed[312],seed[1571],seed[3218],seed[2406],seed[1556],seed[1934],seed[2087],seed[3442],seed[1494],seed[1372],seed[2693],seed[2648],seed[1008],seed[469],seed[2810],seed[3301],seed[2738],seed[3605],seed[3060],seed[2356],seed[1986],seed[2742],seed[1753],seed[2565],seed[344],seed[2522],seed[515],seed[2439],seed[3796],seed[807],seed[3905],seed[547],seed[2197],seed[2947],seed[2656],seed[1466],seed[2544],seed[3578],seed[2746],seed[1327],seed[2647],seed[2140],seed[2335],seed[2194],seed[2906],seed[3898],seed[3689],seed[1687],seed[1508],seed[1801],seed[505],seed[3624],seed[2036],seed[2282],seed[225],seed[1389],seed[1376],seed[1044],seed[1124],seed[1957],seed[1963],seed[1218],seed[1410],seed[1750],seed[149],seed[1330],seed[985],seed[2042],seed[619],seed[3912],seed[1134],seed[3000],seed[876],seed[72],seed[1135],seed[2995],seed[3937],seed[1997],seed[207],seed[1890],seed[1799],seed[2411],seed[1489],seed[329],seed[3660],seed[808],seed[2927],seed[3504],seed[696],seed[1184],seed[320],seed[1949],seed[1666],seed[1294],seed[3351],seed[1848],seed[834],seed[3047],seed[3584],seed[2423],seed[4050],seed[2856],seed[1206],seed[2128],seed[585],seed[2124],seed[3800],seed[3231],seed[795],seed[0],seed[502],seed[41],seed[1590],seed[2495],seed[973],seed[903],seed[126],seed[2387],seed[3230],seed[1194],seed[1593],seed[3748],seed[2878],seed[2498],seed[1718],seed[3402],seed[315],seed[812],seed[3394],seed[4051],seed[3254],seed[2899],seed[1999],seed[1459],seed[1433],seed[2547],seed[3817],seed[2599],seed[2365],seed[2596],seed[2239],seed[3208],seed[940],seed[3372],seed[1420],seed[3387],seed[3343],seed[902],seed[2035],seed[1464],seed[2727],seed[1998],seed[2925],seed[3016],seed[1982],seed[1178],seed[2576],seed[3779],seed[1186],seed[162],seed[2404],seed[3159],seed[3787],seed[1258],seed[2749],seed[2004],seed[3682],seed[1273],seed[442],seed[263],seed[430],seed[2905],seed[38],seed[3226],seed[2066],seed[1960],seed[694],seed[304],seed[1092],seed[3094],seed[951],seed[164],seed[700],seed[1463],seed[1093],seed[1418],seed[2012],seed[797],seed[923],seed[1193],seed[124],seed[20],seed[1262],seed[2354],seed[3073],seed[1020],seed[3596],seed[460],seed[2812],seed[2295],seed[2266],seed[1314],seed[2782],seed[3562],seed[420],seed[949],seed[2388],seed[3495],seed[3176],seed[2473],seed[3552],seed[2014],seed[314],seed[1255],seed[50],seed[2525],seed[1039],seed[529],seed[2722],seed[3758],seed[1926],seed[3297],seed[2465],seed[2790],seed[3821],seed[944],seed[517],seed[1146],seed[2710],seed[28],seed[1277],seed[3431],seed[2122],seed[441],seed[496],seed[2447],seed[3671],seed[3506],seed[2115],seed[1455],seed[1563],seed[2962],seed[1732],seed[3432],seed[3236],seed[519],seed[2921],seed[1985],seed[2930],seed[3847],seed[1891],seed[2459],seed[1574],seed[831],seed[996],seed[3319],seed[1608],seed[991],seed[2653],seed[981],seed[2043],seed[3309],seed[65],seed[3643],seed[2440],seed[1869],seed[3695],seed[3376],seed[2744],seed[3300],seed[3724],seed[3416],seed[1191],seed[1394],seed[3503],seed[712],seed[1269],seed[3425],seed[732],seed[4062],seed[426],seed[2671],seed[2629],seed[1270],seed[776],seed[814],seed[1079],seed[380],seed[2148],seed[2293],seed[2060],seed[3050],seed[1371],seed[2349],seed[4007],seed[2835],seed[2696],seed[2730],seed[3593],seed[3112],seed[2208],seed[2428],seed[2745],seed[3214],seed[2538],seed[3851],seed[1083],seed[1103],seed[1646],seed[676],seed[2956],seed[1402],seed[3813],seed[3433],seed[3401],seed[2130],seed[3240],seed[326],seed[35],seed[2171],seed[247],seed[189],seed[3429],seed[761],seed[1144],seed[2608],seed[1683],seed[4008],seed[2996],seed[555],seed[2971],seed[2517],seed[2773],seed[2959],seed[1847],seed[3579],seed[569],seed[3168],seed[1106],seed[1981],seed[2142],seed[3427],seed[237],seed[1082],seed[2275],seed[1373],seed[287],seed[2928],seed[3520],seed[1030],seed[2747],seed[1930],seed[208],seed[3806],seed[1672],seed[1689],seed[3903],seed[456],seed[1279],seed[1578],seed[1525],seed[3184],seed[2994],seed[3505],seed[3793],seed[1897],seed[1045],seed[1707],seed[1266],seed[122],seed[3901],seed[2924],seed[514],seed[369],seed[3457],seed[3681],seed[2378],seed[3367],seed[378],seed[3305],seed[1915],seed[3085],seed[2564],seed[3325],seed[550],seed[1509],seed[2330],seed[3324],seed[1275],seed[2532],seed[1102],seed[2665],seed[2784],seed[2367],seed[3071],seed[2724],seed[777],seed[4029],seed[2381],seed[1535],seed[953],seed[1132],seed[2602],seed[3939],seed[2200],seed[1638],seed[3914],seed[533],seed[434],seed[3768],seed[2167],seed[3990],seed[165],seed[1645],seed[2352],seed[2676],seed[2658],seed[234],seed[448],seed[258],seed[482],seed[2467],seed[413],seed[4049],seed[2048],seed[3762],seed[2344],seed[2981],seed[2416],seed[538],seed[715],seed[2348],seed[3417],seed[2531],seed[418],seed[3274],seed[589],seed[3861],seed[919],seed[2007],seed[3639],seed[1413],seed[1878],seed[2207],seed[662],seed[790],seed[3488],seed[911],seed[1263],seed[1684],seed[3233],seed[2796],seed[3680],seed[830],seed[1313],seed[2103],seed[2472],seed[3959],seed[1334],seed[2914],seed[1865],seed[1702],seed[3022],seed[2803],seed[1034],seed[242],seed[523],seed[2787],seed[4031],seed[1022],seed[1549],seed[2273],seed[3068],seed[874],seed[2262],seed[1078],seed[274],seed[3776],seed[3672],seed[1853],seed[2876],seed[232],seed[2707],seed[3360],seed[1941],seed[2415],seed[1058],seed[2125],seed[2420],seed[466],seed[146],seed[1029],seed[2751],seed[4040],seed[1828],seed[1174],seed[231],seed[2074],seed[1367],seed[4088],seed[3118],seed[1260],seed[1253],seed[613],seed[167],seed[1583],seed[669],seed[1825],seed[3704],seed[2743],seed[348],seed[3117],seed[183],seed[2603],seed[1631],seed[1910],seed[2307],seed[2366],seed[1267],seed[564],seed[4064],seed[3149],seed[371],seed[2896],seed[2395],seed[2999],seed[1806],seed[900],seed[2019],seed[444],seed[1970],seed[2527],seed[3334],seed[1043],seed[2198],seed[3694],seed[1216],seed[3947],seed[959],seed[1038],seed[762],seed[2988],seed[914],seed[3531],seed[73],seed[4077],seed[1307],seed[404],seed[3705],seed[3641],seed[1150],seed[3933],seed[2316],seed[2637],seed[1182],seed[2355],seed[1567],seed[2497],seed[3970],seed[3586],seed[236],seed[1456],seed[18],seed[1539],seed[3485],seed[2689],seed[2886],seed[3354],seed[3803],seed[2536],seed[2567],seed[3167],seed[638],seed[1800],seed[3467],seed[3113],seed[2687],seed[243],seed[3051],seed[3785],seed[2587],seed[1268],seed[1585],seed[2861],seed[3550],seed[1780],seed[2780],seed[4041],seed[2943],seed[1625],seed[4018],seed[36],seed[3899],seed[2859],seed[3346],seed[660],seed[2890],seed[3981],seed[1049],seed[3538],seed[4026],seed[3955],seed[3210],seed[3675],seed[2068],seed[799],seed[631],seed[2425],seed[431],seed[1765],seed[2860],seed[352],seed[1126],seed[741],seed[2543],seed[1396],seed[259],seed[658],seed[2813],seed[1618],seed[939],seed[1284],seed[63],seed[2686],seed[1077],seed[1002],seed[2049],seed[3067],seed[3368],seed[3272],seed[3311],seed[3713],seed[657],seed[1303],seed[3891],seed[2345],seed[868],seed[2059],seed[2391],seed[4009],seed[2110],seed[859],seed[3994],seed[3189],seed[1874],seed[3373],seed[787],seed[26],seed[1325],seed[3147],seed[1070],seed[3907],seed[3175],seed[3897],seed[1235],seed[1109],seed[1308],seed[3024],seed[1793],seed[3307],seed[1431],seed[863],seed[1783],seed[467],seed[2073],seed[2199],seed[134],seed[2634],seed[1486],seed[257],seed[2086],seed[1880],seed[1151],seed[3090],seed[2146],seed[974],seed[2627],seed[318],seed[3268],seed[2259],seed[3420],seed[3612],seed[791],seed[372],seed[2287],seed[52],seed[1315],seed[268],seed[2136],seed[1072],seed[1110],seed[908],seed[2308],seed[1329],seed[3594],seed[551],seed[144],seed[2703],seed[3095],seed[3227],seed[1318],seed[3143],seed[1434],seed[1054],seed[384],seed[898],seed[1492],seed[3732],seed[3963],seed[196],seed[1770],seed[471],seed[1408],seed[1860],seed[2786],seed[1286],seed[989],seed[3878],seed[3479],seed[1427],seed[2471],seed[2794],seed[600],seed[4061],seed[1570],seed[2119],seed[3743],seed[358],seed[1175],seed[248],seed[2096],seed[2848],seed[3291],seed[2206],seed[1426],seed[1713],seed[1691],seed[3603],seed[2550],seed[1842],seed[3871],seed[3041],seed[748],seed[4055],seed[2433],seed[594],seed[338],seed[2846],seed[636],seed[2549],seed[1771],seed[2523],seed[2179],seed[982],seed[2983],seed[2533],seed[1643],seed[3756],seed[3589],seed[3805],seed[414],seed[3975],seed[1648],seed[1397],seed[1239],seed[3475],seed[1548],seed[796],seed[2247],seed[1024],seed[2407],seed[119],seed[869],seed[2152],seed[3618],seed[2654],seed[2419],seed[689],seed[350],seed[999],seed[3968],seed[2158],seed[2877],seed[1208],seed[3760],seed[3749],seed[2768],seed[3980],seed[3554],seed[120],seed[1749],seed[1742],seed[3169],seed[1591],seed[2977],seed[2177],seed[355],seed[2394],seed[3129],seed[2808],seed[3486],seed[3696],seed[1579],seed[310],seed[1615],seed[3303],seed[2217],seed[3321],seed[449],seed[55],seed[3674],seed[148],seed[2009],seed[2697],seed[2845],seed[2975],seed[552],seed[1248],seed[1497],seed[1010],seed[3223],seed[279],seed[3128],seed[3927],seed[1152],seed[2150],seed[1560],seed[804],seed[3234],seed[3141],seed[2838],seed[1708],seed[2733],seed[157],seed[1907],seed[2958],seed[1623],seed[3322],seed[1789],seed[3708],seed[143],seed[826],seed[1354],seed[336],seed[1526],seed[319],seed[579],seed[850],seed[586],seed[2837],seed[2123],seed[190],seed[107],seed[351],seed[692],seed[1909],seed[3500],seed[6],seed[1296],seed[2559],seed[1820],seed[1942],seed[1052],seed[3876],seed[2098],seed[2143],seed[702],seed[3207],seed[3191],seed[3537],seed[2781],seed[23],seed[1019],seed[2281],seed[2001],seed[1220],seed[610],seed[3881],seed[91],seed[1341],seed[2120],seed[3515],seed[1515],seed[1659],seed[2153],seed[1063],seed[408],seed[4074],seed[3163],seed[1451],seed[3654],seed[3438],seed[3913],seed[3317],seed[2057],seed[1745],seed[3304],seed[1305],seed[2551],seed[971],seed[3638],seed[4067],seed[3684],seed[2731],seed[1348],seed[1725],seed[381],seed[2163],seed[1901],seed[3630],seed[3142],seed[1225],seed[2577],seed[3410],seed[3786],seed[544],seed[1831],seed[291],seed[878],seed[3070],seed[1465],seed[2085],seed[2867],seed[893],seed[1071],seed[665],seed[1792],seed[3172],seed[1617],seed[2225],seed[3610],seed[2759],seed[2623],seed[815],seed[2135],seed[3106],seed[1918],seed[104],seed[391],seed[2521],seed[1719],seed[1232],seed[504],seed[301],seed[948],seed[2232],seed[3145],seed[3996],seed[2181],seed[1927],seed[54],seed[246],seed[3754],seed[3296],seed[2093],seed[4],seed[518],seed[3784],seed[2668],seed[3295],seed[2493],seed[1285],seed[1845],seed[3774],seed[3422],seed[1966],seed[412],seed[2800],seed[1379],seed[2100],seed[402],seed[3253],seed[84],seed[3807],seed[3828],seed[1856],seed[2620],seed[4013],seed[141],seed[2038],seed[3374],seed[2913],seed[1882],seed[848],seed[2636],seed[3493],seed[1490],seed[3017],seed[1699],seed[2319],seed[677],seed[3588],seed[40],seed[3077],seed[2155],seed[2968],seed[3235],seed[705],seed[3508],seed[2005],seed[32],seed[2409],seed[1569],seed[2675],seed[3035],seed[76],seed[1155],seed[2664],seed[1572],seed[3428],seed[1336],seed[4015],seed[1829],seed[1530],seed[2606],seed[1042],seed[2041],seed[857],seed[2540],seed[3739],seed[3855],seed[896],seed[3252],seed[1355],seed[3582],seed[3686],seed[3213],seed[1074],seed[3138],seed[3476],seed[306],seed[2748],seed[309],seed[856],seed[2470],seed[781],seed[3250],seed[2210],seed[535],seed[3962],seed[1064],seed[2823],seed[2323],seed[446],seed[1844],seed[1243],seed[3652],seed[424],seed[1197],seed[1219],seed[3314],seed[2907],seed[531],seed[3201],seed[3444],seed[5],seed[169],seed[864],seed[3964],seed[3440],seed[3809],seed[2053],seed[2075],seed[2218],seed[918],seed[1991],seed[1817],seed[2866],seed[618],seed[1704],seed[1762],seed[2328],seed[4046],seed[1900],seed[3115],seed[1369],seed[763],seed[1236],seed[191],seed[3693],seed[2157],seed[98],seed[2973],seed[1366],seed[2916],seed[102],seed[295],seed[3802],seed[745],seed[3556],seed[2376],seed[1627],seed[2236],seed[2434],seed[174],seed[2510],seed[588],seed[933],seed[3735],seed[1339],seed[998],seed[548],seed[1931],seed[909],seed[1483],seed[798],seed[1224],seed[1240],seed[2254],seed[2405],seed[2195],seed[2901],seed[1794],seed[4072],seed[601],seed[2557],seed[1894],seed[226],seed[1381],seed[1417],seed[1297],seed[2088],seed[1682],seed[1737],seed[616],seed[1936],seed[390],seed[2604],seed[1823],seed[2230],seed[2134],seed[3928],seed[3759],seed[1883],seed[1457],seed[2456],seed[3604],seed[4086],seed[2888],seed[3353],seed[3882],seed[906],seed[3986],seed[3269],seed[1338],seed[3059],seed[1796],seed[766],seed[2505],seed[438],seed[3211],seed[1317],seed[1405],seed[3124],seed[3248],seed[2949],seed[500],seed[2034],seed[3019],seed[1157],seed[3350],seed[1899],seed[363],seed[2340],seed[2723],seed[3012],seed[3767],seed[374],seed[767],seed[2180],seed[3302],seed[2154],seed[3383],seed[2492],seed[1956],seed[3765],seed[2350],seed[1636],seed[1120],seed[2569],seed[1158],seed[3023],seed[2191],seed[3283],seed[1804],seed[428],seed[2201],seed[99],seed[2357],seed[2160],seed[334],seed[595],seed[2220],seed[744],seed[1619],seed[1564],seed[1812],seed[3452],seed[1630],seed[2915],seed[3946],seed[673],seed[1385],seed[34],seed[3798],seed[3263],seed[1575],seed[1710],seed[3645],seed[276],seed[1621],seed[1586],seed[1346],seed[3197],seed[2612],seed[1498],seed[2441],seed[3555],seed[3221],seed[3997],seed[477],seed[4023],seed[541],seed[3323],seed[2375],seed[2639],seed[139],seed[494],seed[2885],seed[293],seed[289],seed[15],seed[308],seed[1416],seed[3080],seed[1430],seed[3615],seed[3518],seed[1040],seed[4016],seed[774],seed[1946],seed[2358],seed[1577],seed[3472],seed[436],seed[3698],seed[2836],seed[2165],seed[706],seed[3753],seed[1965],seed[2410],seed[3243],seed[1055],seed[198],seed[913],seed[1478],seed[2643],seed[2944],seed[419],seed[1411],seed[300],seed[1261],seed[1283],seed[3443],seed[3462],seed[3202],seed[2851],seed[347],seed[345],seed[349],seed[97],seed[3205],seed[938],seed[565],seed[917],seed[3773],seed[3007],seed[3703],seed[439],seed[961],seed[825],seed[2509],seed[634],seed[1211],seed[3870],seed[1641],seed[1399],seed[3661],seed[2284],seed[1179],seed[1650],seed[1700],seed[3078],seed[3193],seed[112],seed[1573],seed[286],seed[1721],seed[3606],seed[3421],seed[2234],seed[546],seed[3460],seed[987],seed[3260],seed[1018],seed[2032],seed[2435],seed[170],seed[986],seed[2235],seed[2552],seed[29],seed[2545],seed[960],seed[3459],seed[755],seed[3087],seed[1495],seed[2222],seed[2605],seed[2421],seed[1594],seed[2468],seed[2080],seed[3716],seed[1872],seed[2186],seed[1557],seed[2788],seed[2933],seed[1068],seed[4035],seed[3312],seed[3086],seed[1724],seed[1599],seed[2306],seed[2214],seed[2777],seed[3228],seed[4038],seed[3458],seed[1123],seed[1095],seed[1596],seed[3795],seed[1364],seed[2487],seed[187],seed[1972],seed[2558],seed[711],seed[1470],seed[3829],seed[3764],seed[2957],seed[1080],seed[1923],seed[1589],seed[3804],seed[324],seed[3185],seed[3718],seed[95],seed[1868],seed[2107],seed[1419],seed[1674],seed[1300],seed[1004],seed[1581],seed[3101],seed[839],seed[2990],seed[653],seed[645],seed[3182],seed[3761],seed[2572],seed[3585],seed[3229],seed[3042],seed[3527],seed[1108],seed[1983],seed[3904],seed[823],seed[2582],seed[1013],seed[3238],seed[137],seed[1065],seed[2919],seed[2900],seed[1037],seed[2613],seed[1370],seed[2283],seed[3885],seed[1447],seed[3399],seed[39],seed[1864],seed[2678],seed[3146],seed[1522],seed[2017],seed[3406],seed[415],seed[1808],seed[2633],seed[3583],seed[967],seed[2984],seed[643],seed[3183],seed[480],seed[1827],seed[184],seed[2322],seed[521],seed[786],seed[166],seed[2698],seed[1171],seed[1047],seed[140],seed[806],seed[3571],seed[3580],seed[3563],seed[867],seed[822],seed[805],seed[3621],seed[445],seed[94],seed[3247],seed[1814],seed[4048],seed[2511],seed[553],seed[1747],seed[1566],seed[2708],seed[604],seed[719],seed[281],seed[2039],seed[3649],seed[743],seed[3608],seed[96],seed[1006],seed[3382],seed[955],seed[2942],seed[1221],seed[3572],seed[3329],seed[664],seed[1228],seed[2452],seed[3846],seed[979],seed[3179],seed[3364],seed[3573],seed[2716],seed[637],seed[3415],seed[3110],seed[3426],seed[1350],seed[2528],seed[2127],seed[1775],seed[513],seed[2955],seed[1295],seed[2315],seed[1136],seed[3651],seed[599],seed[333],seed[2460],seed[3512],seed[3944],seed[266],seed[2062],seed[1785],seed[3551],seed[3136],seed[3547],seed[739],seed[1154],seed[1819],seed[3858],seed[1395],seed[2249],seed[3430],seed[2018],seed[3498],seed[537],seed[343],seed[2455],seed[110],seed[3257],seed[1507],seed[752],seed[1223],seed[283],seed[3386],seed[570],seed[3046],seed[1094],seed[113],seed[2610],seed[48],seed[3036],seed[1097],seed[4081],seed[1779],seed[219],seed[159],seed[709],seed[614],seed[197],seed[3950],seed[459],seed[2513],seed[1436],seed[1125],seed[2399],seed[3447],seed[3843],seed[782],seed[4093],seed[3519],seed[3490],seed[688],seed[925],seed[2820],seed[296],seed[3564],seed[3734],seed[3126],seed[1656],seed[1818],seed[731],seed[1948],seed[2373],seed[215],seed[3745],seed[1473],seed[1101],seed[1562],seed[2109],seed[282],seed[393],seed[540],seed[127],seed[2446],seed[695],seed[305],seed[179],seed[3513],seed[4094],seed[2614],seed[956],seed[770],seed[707],seed[2868],seed[3032],seed[71],seed[227],seed[3670],seed[4039],seed[3987],seed[1458],seed[1384],seed[2638],seed[1335],seed[1375],seed[1086],seed[922],seed[2083],seed[980],seed[4014],seed[847],seed[1130],seed[727],seed[2518],seed[1160],seed[560],seed[682],seed[2324],seed[2641],seed[2674],seed[3043],seed[202],seed[3190],seed[3867],seed[3181],seed[2161],seed[3546],seed[3710],seed[524],seed[2556],seed[57],seed[322],seed[621],seed[687],seed[152],seed[2454],seed[532],seed[2884],seed[405],seed[3967],seed[2524],seed[3216],seed[2116],seed[2726],seed[2824],seed[3511],seed[3799],seed[2337],seed[1438],seed[697],seed[2298],seed[3626],seed[3166],seed[1993],seed[2893],seed[1944],seed[1746],seed[88],seed[3326],seed[3533],seed[3791],seed[203],seed[1639],seed[3403],seed[3771],seed[2078],seed[2385],seed[907],seed[3741],seed[1634],seed[603],seed[1561],seed[3892],seed[3909],seed[2684],seed[2765],seed[2309],seed[3900],seed[3966],seed[3969],seed[904],seed[2445],seed[3516],seed[2095],seed[2855],seed[370],seed[273],seed[69],seed[3008],seed[627],seed[1678],seed[58],seed[3424],seed[3816],seed[1272],seed[3053],seed[3196],seed[3448],seed[1609],seed[800],seed[4075],seed[37],seed[2546],seed[2147],seed[2611],seed[2169],seed[2669],seed[3011],seed[3542],seed[2826],seed[2226],seed[3337],seed[1181],seed[2579],seed[2246],seed[1958],seed[3108],seed[3535],seed[1604],seed[3148],seed[1802],seed[587],seed[3747],seed[406],seed[2029],seed[396],seed[3917],seed[1359],seed[1140],seed[1772],seed[2327],seed[2002],seed[2898],seed[932],seed[4092],seed[2805],seed[1099],seed[3543],seed[3310],seed[3971],seed[1041],seed[1007],seed[1688],seed[2263],seed[788],seed[2216],seed[1654],seed[1050],seed[1754],seed[1813],seed[3926],seed[757],seed[16],seed[3015],seed[1889],seed[4070],seed[2535],seed[3418],seed[2767],seed[2368],seed[720],seed[3481],seed[2461],seed[2624],seed[644],seed[3951],seed[353],seed[3276],seed[3203],seed[1111],seed[954],seed[1588],seed[2750],seed[849],seed[155],seed[1787],seed[3290],seed[3920],seed[773],seed[886],seed[2408],seed[4000],seed[2000],seed[1544],seed[1720],seed[1782],seed[394],seed[3125],seed[3135],seed[2929],seed[1028],seed[2849],seed[3150],seed[2432],seed[680],seed[1803],seed[3812],seed[646],seed[3133],seed[465],seed[3206],seed[3976],seed[3392],seed[3685],seed[1658],seed[3152],seed[316],seed[117],seed[765],seed[3120],seed[1301],seed[2051],seed[2390],seed[1343],seed[3865],seed[725],seed[635],seed[3746],seed[3781],seed[1360],seed[2632],seed[2317],seed[2954],seed[3541],seed[591],seed[3888],seed[1026],seed[2903],seed[3278],seed[3737],seed[1199],seed[3497],seed[1468],seed[1693],seed[2046],seed[2227],seed[2706],seed[1250],seed[175],seed[4005],seed[2334],seed[3834],seed[136],seed[3841],seed[3666],seed[3161],seed[4024],seed[45],seed[3173],seed[2371],seed[1928],seed[947],seed[2574],seed[2052],seed[1711],seed[2065],seed[1462],seed[25],seed[1809],seed[3908],seed[2694],seed[3001],seed[3154],seed[2187],seed[1886],seed[368],seed[70],seed[2037],seed[2869],seed[659],seed[1059],seed[1955],seed[2772],seed[1729],seed[1922],seed[462],seed[180],seed[3013],seed[79],seed[3688],seed[2619],seed[3923],seed[1962],seed[3127],seed[2449],seed[2300],seed[3464],seed[2829],seed[3995],seed[3998],seed[1546],seed[3251],seed[331],seed[2500],seed[1051],seed[3780],seed[2850],seed[2508],seed[2704],seed[1119],seed[3832],seed[3111],seed[3823],seed[1551],seed[261],seed[86],seed[2402],seed[3249],seed[2600],seed[2031],seed[3599],seed[1163],seed[995],seed[1264],seed[506],seed[1309],seed[3171],seed[1472],seed[1776],seed[2104],seed[2753],seed[2437],seed[2666],seed[2296],seed[130],seed[2774],seed[2809],seed[1622],seed[3316],seed[1502],seed[1057],seed[1857],seed[172],seed[2677],seed[3974],seed[835],seed[3186],seed[1690],seed[3931],seed[789],seed[1159],seed[12],seed[2681],seed[2909],seed[2662],seed[2622],seed[1837],seed[2172],seed[2895],seed[1252],seed[2737],seed[3943],seed[1714],seed[2961],seed[3544],seed[3863],seed[3393],seed[3217],seed[1241],seed[1815],seed[3062],seed[2013],seed[654],seed[2691],seed[3066],seed[3455],seed[1701],seed[1345],seed[31],seed[3930],seed[2325],seed[89],seed[1835],seed[2872],seed[3553],seed[488],seed[1517],seed[3461],seed[2444],seed[3239],seed[2649],seed[509],seed[2336],seed[2310],seed[373],seed[2431],seed[1696],seed[2739],seed[3751],seed[2418],seed[3277],seed[461],seed[3906],seed[2276],seed[3866],seed[3451],seed[1293],seed[2070],seed[3242],seed[173],seed[1512],seed[1249],seed[1524],seed[3794],seed[3099],seed[683],seed[2858],seed[733],seed[1227],seed[3646],seed[417],seed[1011],seed[3857],seed[3524],seed[670],seed[103],seed[2028],seed[4030],seed[407],seed[574],seed[46],seed[2190],seed[2979],seed[819],seed[290],seed[2997],seed[4032],seed[1190],seed[1832],seed[3595],seed[195],seed[3935],seed[821],seed[978],seed[83],seed[2166],seed[1195],seed[3956],seed[2185],seed[2079],seed[3522],seed[704],seed[142],seed[615],seed[1187],seed[1892],seed[2286],seed[2288],seed[3140],seed[1009],seed[1734],seed[3289],seed[47],seed[816],seed[1319],seed[3293],seed[3348],seed[366],seed[400],seed[2364],seed[3709],seed[1117],seed[1774],seed[210],seed[1821],seed[2950],seed[1424],seed[2804],seed[2091],seed[185],seed[44],seed[342],seed[129],seed[1316],seed[3003],seed[3782],seed[1628],seed[2761],seed[3830],seed[3049],seed[3371],seed[3984],seed[1387],seed[2617],seed[539],seed[1705],seed[49],seed[3788],seed[2010],seed[2040],seed[1204],seed[3355],seed[2429],seed[794],seed[3752],seed[3407],seed[1302],seed[1471],seed[2277],seed[199],seed[171],seed[1292],seed[1651],seed[1558],seed[1475],seed[2030],seed[3662],seed[3338],seed[916],seed[3778],seed[1398],seed[2114],seed[935],seed[3730],seed[1185],seed[675],seed[2099],seed[397],seed[272],seed[1552],seed[2542],seed[2779],seed[3985],seed[582],seed[2891],seed[2635],seed[2519],seed[3031],seed[2274],seed[440],seed[581],seed[2285],seed[3558],seed[703],seed[1924],seed[1153],seed[2626],seed[921],seed[1968],seed[2121],seed[2789],seed[2174],seed[3419],seed[1875],seed[327],seed[317],seed[3391],seed[2601],seed[3978],seed[802],seed[1365],seed[912],seed[2887],seed[4037],seed[3330],seed[2964],seed[1450],seed[377],seed[220],seed[1021],seed[1511],seed[3105],seed[3992],seed[3219],seed[2486],seed[1602],seed[1353],seed[128],seed[4006],seed[1349],seed[2178],seed[325],seed[642],seed[678],seed[690],seed[3332],seed[11],seed[454],seed[1740],seed[3076],seed[716],seed[629],seed[2205],seed[3561],seed[3294],seed[1382],seed[161],seed[3559],seed[1180],seed[153],seed[1769],seed[1344],seed[367],seed[1743],seed[3972],seed[2770],seed[43],seed[1598],seed[339],seed[571],seed[2864],seed[1554],seed[557],seed[1597],seed[1129],seed[1445],seed[1407],seed[3845],seed[2948],seed[1662],seed[1453],seed[3162],seed[3093],seed[1166],seed[2311],seed[2250],seed[1242],seed[93],seed[475],seed[2261],seed[292],seed[803],seed[255],seed[4002],seed[2875],seed[2660],seed[1107],seed[1217],seed[2575],seed[2935],seed[3040],seed[2025],seed[3854],seed[1735],seed[2360],seed[829],seed[229],seed[1781],seed[3844],seed[1854],seed[2963],seed[7],seed[1031],seed[699],seed[1491],seed[993],seed[846],seed[211],seed[87],seed[1352],seed[1777],seed[3299],seed[205],seed[2329],seed[2515],seed[734],seed[1679],seed[2491],seed[3137],seed[2221],seed[3648],seed[3569],seed[132],seed[3530],seed[2873],seed[1056],seed[3098],seed[2842],seed[3097],seed[3570],seed[768],seed[1192],seed[742],seed[2370],seed[1974],seed[3204],seed[2966],seed[158],seed[1971],seed[1333],seed[1061],seed[647],seed[2897],seed[3625],seed[2458],seed[297],seed[3665],seed[1992],seed[2346],seed[3942],seed[738],seed[3489],seed[2987],seed[2347],seed[1276],seed[3441],seed[1778],seed[3676],seed[495],seed[545],seed[3083],seed[1046],seed[2917],seed[254],seed[2457],seed[968],seed[1500],seed[889],seed[997],seed[556],seed[1053],seed[2507],seed[606],seed[2553],seed[2450],seed[3390],seed[3818],seed[785],seed[2688],seed[3057],seed[3212],seed[1712],seed[1885],seed[962],seed[4034],seed[2326],seed[3777],seed[3039],seed[975],seed[2938],seed[2240],seed[3770],seed[2237],seed[2985],seed[2430],seed[3678],seed[3096],seed[2003],seed[2170],seed[357],seed[3054],seed[2644],seed[1840],seed[2453],seed[3723],seed[3952],seed[3576],seed[2481],seed[4063],seed[1446],seed[1532],seed[1210],seed[2314],seed[3139],seed[303],seed[2269],seed[1984],seed[1168],seed[62],seed[403],seed[1506],seed[3839],seed[2202],seed[717],seed[3144],seed[4065],seed[1685],seed[1320],seed[1670],seed[2392],seed[3958],seed[3158],seed[1811],seed[860],seed[3957],seed[2268],seed[13],seed[133],seed[3104],seed[686],seed[3915],seed[222],seed[3597],seed[2778],seed[2094],seed[853],seed[213],seed[977],seed[3091],seed[708],seed[3496],seed[1245],seed[3528],seed[758],seed[3617],seed[2252],seed[1726],seed[1518],seed[3640],seed[2760],seed[4079],seed[3581],seed[3815],seed[3450],seed[8],seed[1172],seed[468],seed[976],seed[1988],seed[1298],seed[1994],seed[498],seed[332],seed[3408],seed[1866],seed[879],seed[90],seed[3288],seed[2506],seed[1452],seed[1404],seed[1257],seed[3514],seed[2442],seed[2970],seed[861],seed[2182],seed[1202],seed[2379],seed[64],seed[1605],seed[2892],seed[596],seed[840],seed[592],seed[520],seed[1969],seed[651],seed[3949],seed[3187],seed[3255],seed[899],seed[399],seed[2673],seed[1282],seed[1541],seed[1147],seed[630],seed[1176],seed[2102],seed[115],seed[1089],seed[1493],seed[1680],seed[3766],seed[1805],seed[2798],seed[1441],seed[2802],seed[3331],seed[2562],seed[256],seed[1016],seed[3993],seed[3306],seed[942],seed[3921],seed[2797],seed[3339],seed[931],seed[2874],seed[100],seed[3044],seed[684],seed[2862],seed[1036],seed[2854],seed[1616],seed[2571],seed[2297],seed[3653],seed[929],seed[3848],seed[3954],seed[302],seed[2597],seed[1917],seed[2537],seed[1728],seed[275],seed[249],seed[2264],seed[575],seed[723],seed[463],seed[1014],seed[1613],seed[844],seed[1290],seed[1278],seed[756],seed[2847],seed[1698],seed[2819],seed[3484],seed[188],seed[59],seed[623],seed[3079],seed[3862],seed[2936],seed[1480],seed[2301],seed[3285],seed[2072],seed[244],seed[3690],seed[984],seed[3010],seed[2616],seed[1066],seed[722],seed[3357],seed[1836],seed[453],seed[3824],seed[1337],seed[2257],seed[928],seed[3894],seed[3775],seed[1164],seed[2006],seed[1281],seed[1768],seed[3412],seed[3929],seed[3801],seed[2714],seed[1306],seed[2700],seed[3864],seed[1487],seed[2563],seed[3258],seed[1391],seed[2870],seed[3902],seed[1076],seed[779],seed[125],seed[554],seed[2960],seed[1881],seed[666],seed[1989],seed[2830],seed[945],seed[455],seed[2490],seed[988],seed[2480],seed[2712],seed[2766],seed[1888],seed[1448],seed[3790],seed[2554],seed[1862],seed[2464],seed[437],seed[609],seed[1128],seed[2776],seed[1861],seed[3072],seed[941],seed[2530],seed[2534],seed[837],seed[1741],seed[910],seed[1527],seed[648],seed[3377],seed[299],seed[1386],seed[663],seed[395],seed[2682],seed[3711],seed[2426],seed[1331],seed[4010],seed[108],seed[3808],seed[2692],seed[3232],seed[3634],seed[625],seed[1167],seed[1607],seed[3849],seed[3601],seed[2241],seed[1173],seed[3609],seed[1786],seed[3164],seed[2145],seed[3627],seed[398],seed[3655],seed[3600],seed[2231],seed[3423],seed[2332],seed[3246],seed[969],seed[1833],seed[1788],seed[1012],seed[239],seed[401],seed[3567],seed[1113],seed[843],seed[583],seed[926],seed[1576],seed[3463],seed[1025],seed[1987],seed[3414],seed[3629],seed[2670],seed[875],seed[3814],seed[4090],seed[2756],seed[1],seed[2585],seed[3717],seed[2427],seed[3523],seed[2389],seed[572],seed[2646],seed[2292],seed[2338],seed[238],seed[217],seed[2578],seed[4019],seed[877],seed[512],seed[1841],seed[1846],seed[2588],seed[1933],seed[965],seed[2401],seed[1790],seed[156],seed[1085],seed[3132],seed[2016],seed[486],seed[2484],seed[1816],seed[2713],seed[510],seed[427],seed[3284],seed[2980],seed[2496],seed[3568],seed[3029],seed[1896],seed[1996],seed[2541],seed[972],seed[2438],seed[1400],seed[3560],seed[1356],seed[1759],seed[801],seed[2520],seed[3591],seed[3647],seed[3473],seed[2952],seed[679],seed[2566],seed[1481],seed[3400],seed[892],seed[2881],seed[2020],seed[3874],seed[1555],seed[1727],seed[77],seed[1401],seed[193],seed[3347],seed[3669],seed[4020],seed[201],seed[1488],seed[2672],seed[1460],seed[668],seed[3619],seed[534],seed[598],seed[3177],seed[602],seed[1751],seed[1839],seed[718],seed[3273],seed[2699],seed[1758],seed[2655],seed[1437],seed[2642],seed[2258],seed[2118],seed[2412],seed[288],seed[4036],seed[890],seed[3611],seed[1288],seed[4047],seed[1838],seed[3840],seed[3499],seed[2941],seed[1547],seed[1947],seed[1482],seed[597],seed[147],seed[2501],seed[2063],seed[3075],seed[3719],seed[3507],seed[2799],seed[1048],seed[154],seed[842],seed[2290],seed[3733],seed[754],seed[3534],seed[2203],seed[970],seed[3953],seed[364],seed[307],seed[501],seed[3859],seed[2248],seed[4057],seed[3725],seed[2398],seed[1467],seed[269],seed[3081],seed[1403],seed[186],seed[2448],seed[176],seed[432],seed[2047],seed[3936],seed[2793],seed[836],seed[1767],seed[824],seed[2573],seed[1697],seed[1870],seed[966],seed[233],seed[375],seed[423],seed[2735],seed[1528],seed[2215],seed[2911],seed[2092],seed[661],seed[1358],seed[1138],seed[3379],seed[2343],seed[150],seed[2108],seed[429],seed[386],seed[2469],seed[2806],seed[3736],seed[671],seed[1069],seed[3650],seed[1000],seed[1501],seed[3783],seed[2024],seed[3509],seed[1311],seed[2112],seed[1671],seed[433],seed[123],seed[2305],seed[1504],seed[3385],seed[3396],seed[710],seed[2920],seed[2992],seed[3397],seed[3721],seed[2238],seed[1663],seed[891],seed[2514],seed[3982],seed[2397],seed[2974],seed[335],seed[1752],seed[3027],seed[3707],seed[2512],seed[2244],seed[2321],seed[2245],seed[2640],seed[628],seed[2932],seed[2333],seed[4033],seed[1629],seed[3266],seed[881],seed[497],seed[3769],seed[2113],seed[4058],seed[730],seed[2105],seed[1521],seed[3973],seed[3114],seed[3940],seed[1499],seed[3644],seed[3267],seed[3109],seed[1939],seed[3292],seed[387],seed[51],seed[2539],seed[3056],seed[3979],seed[612],seed[2228],seed[746],seed[3103],seed[3545],seed[3313],seed[2757],seed[3262],seed[75],seed[2822],seed[3005],seed[4066],seed[221],seed[721],seed[1112],seed[385],seed[769],seed[1357],seed[530],seed[493],seed[1640],seed[3123],seed[3510],seed[2097],seed[2982],seed[3404],seed[2607],seed[2383],seed[3026],seed[3557],seed[1736],seed[3726],seed[2377],seed[992],seed[735],seed[1748],seed[3880],seed[1925],seed[2156],seed[3456],seed[3089],seed[2594],seed[652],seed[2721],seed[1953],seed[1514],seed[2695],seed[2719],seed[2593],seed[3082],seed[1667],seed[2417],seed[3287],seed[3875],seed[1332],seed[2843],seed[1289],seed[1990],seed[1973],seed[1920],seed[845],seed[1657],seed[2910],seed[1945],seed[2618],seed[2403],seed[435],seed[3700],seed[566],seed[1677],seed[1709],seed[1392],seed[792],seed[2595],seed[2631],seed[204],seed[1592],seed[3130],seed[1201],seed[2926],seed[3160],seed[182],seed[4025],seed[1121],seed[2061],seed[3789],seed[3004],seed[1686],seed[450],seed[1200],seed[3637],seed[2785],seed[340],seed[3025],seed[1676],seed[1247],seed[1959],seed[3827],seed[3884],seed[2548],seed[2106],seed[1265],seed[1443],seed[2451],seed[228],seed[42],seed[2705],seed[3058],seed[3668],seed[3856],seed[3501],seed[1203],seed[2840],seed[27],seed[2271],seed[827],seed[1545],seed[525],seed[2598],seed[2922],seed[1660],seed[1023],seed[865],seed[3134],seed[209],seed[2560],seed[3014],seed[346],seed[3633],seed[3587],seed[1921],seed[1764],seed[641],seed[3879],seed[2683],seed[1409],seed[3131],seed[3409],seed[2082],seed[3349],seed[1673],seed[1887],seed[2318],seed[2175],seed[251],seed[3860],seed[1543],seed[379],seed[1444],seed[3195],seed[1580],seed[2775],seed[2055],seed[3842],seed[1624],seed[2151],seed[2242],seed[313],seed[1600],seed[936],seed[894],seed[3642],seed[250],seed[852],seed[200],seed[3318],seed[2734],seed[2144],seed[3437],seed[1474],seed[2320],seed[2953],seed[833],seed[2436],seed[2801],seed[1137],seed[818],seed[905],seed[56],seed[2902],seed[1383],seed[443],seed[3889],seed[3887],seed[2413],seed[2504],seed[1716],seed[1362],seed[2090],seed[1131],seed[3566],seed[1496],seed[1903],seed[2213],seed[2117],seed[280],seed[952],seed[1873],seed[3315],seed[3614],seed[2341],seed[3333],seed[323],seed[1824],seed[3107],seed[2879],seed[2362],seed[2581],seed[2732],seed[3831],seed[2189],seed[2880],seed[1145],seed[1858],seed[2064],seed[2833],seed[2736],seed[1961],seed[4071],seed[1406],seed[2702],seed[298],seed[2584],seed[2393],seed[491],seed[1603],seed[2939],seed[1916],seed[3910],seed[1104],seed[2807],seed[3999],seed[3055],seed[624],seed[543],seed[750],seed[1906],seed[1189],seed[2993],seed[2084],seed[1237],seed[2351],seed[3632],seed[2967],seed[1898],seed[2372],seed[264],seed[2304],seed[3446],seed[2168],seed[1428],seed[2628],seed[2056],seed[3395],seed[3192],seed[964],seed[1516],seed[2589],seed[3549],seed[1717],seed[3256],seed[3712],seed[1479],seed[866],seed[3298],seed[356],seed[1523],seed[2008],seed[360],seed[1584],seed[862],seed[1230],seed[2229],seed[235],seed[206],seed[2853],seed[2353],seed[3453],seed[4054],seed[3465],seed[2591],seed[1188],seed[3853],seed[3502],seed[3590],seed[1170],seed[1234],seed[1952],seed[1538],seed[527],seed[478],seed[2243],seed[3122],seed[729],seed[1649],seed[3835],seed[4089],seed[3362],seed[2791],seed[1723],seed[354],seed[640],seed[3699],seed[2889],seed[3328],seed[194],seed[3714],seed[1027],seed[2289],seed[590],seed[3454],seed[30],seed[1978],seed[1559],seed[3270],seed[21],seed[2081],seed[1116],seed[3153],seed[656],seed[605],seed[1141],seed[1148],seed[1127],seed[177],seed[2821],seed[728],seed[2841],seed[2894],seed[2969],seed[4045],seed[3064],seed[3170],seed[1851],seed[1975],seed[622],seed[3468],seed[3988],seed[2485],seed[212],seed[2192],seed[4056],seed[3245],seed[2044],seed[3100],seed[2679],seed[3281],seed[1035],seed[2054],seed[2568],seed[1156],seed[4004],seed[3225],seed[1100],seed[3540],seed[1606],seed[1142],seed[1757],seed[3358],seed[1212],seed[1761],seed[2312],seed[330],seed[3941],seed[3359],seed[4060],seed[3033],seed[751],seed[473],seed[3602],seed[111],seed[1612],seed[943],seed[1033],seed[3405],seed[3945],seed[3340],seed[2857],seed[883],seed[1280],seed[3613],seed[3525],seed[474],seed[639],seed[780],seed[2022],seed[691],seed[713],seed[3607],seed[3592],seed[1849],seed[2718],seed[1461],seed[2690],seed[1668],seed[511],seed[3469],seed[178],seed[3715],seed[1231],seed[1347],seed[1291],seed[813],seed[3792],seed[311],seed[2752],seed[3002],seed[793],seed[3720],seed[3521],seed[3492],seed[3822],seed[3065],seed[1661],seed[1810],seed[3833],seed[3873],seed[2972],seed[3275],seed[3656],seed[901],seed[2828],seed[3020],seed[2302],seed[3048],seed[3435],seed[4027],seed[3483],seed[138],seed[608],seed[617],seed[2965],seed[3209],seed[2380],seed[1177],seed[1807],seed[4091],seed[2918],seed[2466],seed[3494],seed[884],seed[1198],seed[1937],seed[14],seed[3411],seed[3691],seed[3526],seed[4087],seed[1312],seed[109],seed[1115],seed[1422],seed[1328],seed[1733],seed[421],seed[2609],seed[1852],seed[3006],seed[2462],seed[1763],seed[216],seed[61],seed[2021],seed[1542],seed[82],seed[2923],seed[2253],seed[1477],seed[337],seed[3102],seed[858],seed[2382],seed[1476],seed[1863],seed[1665],seed[576],seed[2291],seed[3342],seed[2313],seed[1871],seed[3045],seed[855],seed[1550],seed[2818],seed[3157],seed[267],seed[3628],seed[3838],seed[1715],seed[3180],seed[508],seed[2255],seed[3308]};
//        seed10 <= {seed[3624],seed[2102],seed[1027],seed[2471],seed[3952],seed[3977],seed[2390],seed[521],seed[611],seed[1731],seed[624],seed[2913],seed[990],seed[1577],seed[3172],seed[80],seed[3010],seed[2263],seed[793],seed[582],seed[2671],seed[3186],seed[1654],seed[2864],seed[199],seed[3321],seed[1964],seed[3311],seed[1230],seed[4060],seed[1850],seed[3641],seed[2979],seed[2823],seed[1375],seed[4041],seed[699],seed[3877],seed[1942],seed[2009],seed[3599],seed[457],seed[1921],seed[3659],seed[2425],seed[3963],seed[2162],seed[861],seed[2616],seed[2987],seed[3047],seed[2444],seed[3861],seed[325],seed[2833],seed[3203],seed[2954],seed[671],seed[1005],seed[2686],seed[112],seed[2034],seed[1420],seed[753],seed[3388],seed[1327],seed[89],seed[202],seed[777],seed[1208],seed[2882],seed[4065],seed[353],seed[2972],seed[1885],seed[190],seed[3],seed[3727],seed[1744],seed[1745],seed[885],seed[77],seed[1185],seed[1038],seed[2600],seed[887],seed[2801],seed[3718],seed[3444],seed[2218],seed[529],seed[680],seed[1879],seed[4066],seed[967],seed[3291],seed[40],seed[3192],seed[3643],seed[238],seed[2769],seed[2052],seed[2473],seed[1514],seed[1310],seed[2347],seed[3269],seed[1968],seed[2876],seed[2412],seed[1549],seed[2664],seed[1379],seed[3839],seed[808],seed[2803],seed[2003],seed[2295],seed[1993],seed[1155],seed[550],seed[700],seed[1334],seed[3306],seed[3316],seed[1153],seed[1837],seed[2525],seed[713],seed[2441],seed[1352],seed[729],seed[64],seed[348],seed[1887],seed[2970],seed[595],seed[3805],seed[1688],seed[870],seed[1233],seed[1878],seed[368],seed[3993],seed[419],seed[4074],seed[274],seed[2279],seed[1930],seed[3268],seed[203],seed[2842],seed[3240],seed[1010],seed[1068],seed[2812],seed[2495],seed[1637],seed[2649],seed[1796],seed[3767],seed[2507],seed[1540],seed[3348],seed[590],seed[2024],seed[3602],seed[50],seed[3353],seed[1762],seed[1965],seed[2221],seed[2054],seed[342],seed[3800],seed[207],seed[2593],seed[1316],seed[3809],seed[1623],seed[6],seed[286],seed[344],seed[2381],seed[3079],seed[1210],seed[2017],seed[1291],seed[302],seed[1363],seed[946],seed[1950],seed[3214],seed[2504],seed[4087],seed[1618],seed[2108],seed[3420],seed[997],seed[371],seed[1365],seed[2258],seed[2070],seed[2701],seed[952],seed[129],seed[2008],seed[3006],seed[16],seed[244],seed[1324],seed[553],seed[3096],seed[367],seed[2318],seed[2532],seed[1227],seed[3329],seed[2627],seed[1404],seed[3971],seed[1614],seed[4059],seed[1458],seed[685],seed[375],seed[3464],seed[1919],seed[2125],seed[2084],seed[773],seed[3666],seed[3127],seed[597],seed[2016],seed[575],seed[1653],seed[1364],seed[1643],seed[489],seed[3499],seed[1106],seed[642],seed[1561],seed[1438],seed[470],seed[18],seed[1289],seed[733],seed[1518],seed[2528],seed[97],seed[544],seed[663],seed[3537],seed[4075],seed[669],seed[1882],seed[3675],seed[3867],seed[888],seed[3872],seed[1550],seed[2937],seed[2784],seed[2486],seed[219],seed[2524],seed[641],seed[31],seed[113],seed[3454],seed[2587],seed[1719],seed[1773],seed[2406],seed[3121],seed[963],seed[1441],seed[973],seed[2091],seed[3290],seed[3275],seed[235],seed[2929],seed[3583],seed[3597],seed[100],seed[2834],seed[3563],seed[2130],seed[2362],seed[2297],seed[2619],seed[1860],seed[3983],seed[2517],seed[3086],seed[467],seed[288],seed[1865],seed[4002],seed[3802],seed[2632],seed[2777],seed[155],seed[3526],seed[3038],seed[622],seed[2299],seed[762],seed[2974],seed[532],seed[1689],seed[1813],seed[410],seed[2774],seed[2867],seed[2621],seed[159],seed[3202],seed[1279],seed[2339],seed[3961],seed[1533],seed[3535],seed[1362],seed[229],seed[1013],seed[4022],seed[554],seed[2180],seed[1666],seed[1682],seed[95],seed[2199],seed[991],seed[123],seed[989],seed[1201],seed[676],seed[471],seed[56],seed[662],seed[3950],seed[1408],seed[1048],seed[1202],seed[29],seed[2531],seed[3881],seed[2661],seed[1353],seed[2436],seed[1923],seed[3387],seed[2958],seed[3527],seed[2626],seed[1121],seed[3441],seed[3572],seed[1248],seed[2107],seed[2004],seed[1803],seed[3377],seed[795],seed[2453],seed[4037],seed[2167],seed[2551],seed[605],seed[694],seed[1394],seed[3492],seed[2676],seed[2918],seed[1284],seed[1736],seed[2432],seed[3631],seed[1576],seed[1782],seed[679],seed[1189],seed[2113],seed[2442],seed[42],seed[486],seed[3895],seed[668],seed[2350],seed[3391],seed[376],seed[2560],seed[1077],seed[2602],seed[1494],seed[3813],seed[1465],seed[426],seed[3147],seed[2206],seed[4025],seed[3264],seed[2492],seed[3518],seed[717],seed[591],seed[2811],seed[160],seed[3515],seed[3789],seed[3978],seed[2591],seed[3610],seed[2831],seed[3236],seed[53],seed[407],seed[381],seed[339],seed[301],seed[3178],seed[953],seed[839],seed[90],seed[1396],seed[3762],seed[3663],seed[2853],seed[581],seed[1370],seed[552],seed[1390],seed[1181],seed[3614],seed[4033],seed[1239],seed[2150],seed[2076],seed[1672],seed[1466],seed[3893],seed[828],seed[2756],seed[2706],seed[652],seed[646],seed[2251],seed[1815],seed[1109],seed[3764],seed[2051],seed[2730],seed[3029],seed[3892],seed[1099],seed[1145],seed[38],seed[2977],seed[718],seed[2982],seed[3953],seed[1501],seed[1816],seed[1806],seed[4034],seed[2061],seed[3104],seed[7],seed[386],seed[2173],seed[8],seed[945],seed[3401],seed[2553],seed[3714],seed[1909],seed[838],seed[1776],seed[3976],seed[3871],seed[2338],seed[3836],seed[1510],seed[1044],seed[2767],seed[1366],seed[3386],seed[380],seed[1030],seed[1384],seed[720],seed[3513],seed[485],seed[3141],seed[3865],seed[3123],seed[2343],seed[3365],seed[2422],seed[2168],seed[2097],seed[2681],seed[2566],seed[3347],seed[3342],seed[304],seed[2576],seed[3571],seed[922],seed[1599],seed[3003],seed[2790],seed[3285],seed[3379],seed[1344],seed[3848],seed[2736],seed[2185],seed[1624],seed[2021],seed[2922],seed[3191],seed[834],seed[1183],seed[3668],seed[2376],seed[2465],seed[1073],seed[3734],seed[3399],seed[1972],seed[3937],seed[975],seed[1276],seed[2253],seed[243],seed[3901],seed[4070],seed[1251],seed[2967],seed[3238],seed[3355],seed[960],seed[4010],seed[142],seed[3906],seed[1931],seed[4067],seed[2928],seed[2691],seed[3065],seed[3448],seed[3325],seed[3590],seed[1246],seed[763],seed[1405],seed[3760],seed[3022],seed[1409],seed[3478],seed[2100],seed[3676],seed[1461],seed[523],seed[463],seed[1709],seed[2605],seed[2244],seed[3480],seed[1794],seed[2692],seed[1301],seed[464],seed[647],seed[545],seed[1308],seed[3930],seed[2386],seed[4021],seed[101],seed[1900],seed[3181],seed[1977],seed[2699],seed[3260],seed[1026],seed[1385],seed[1329],seed[3049],seed[3462],seed[1095],seed[2788],seed[2696],seed[1676],seed[623],seed[1870],seed[2521],seed[3905],seed[854],seed[213],seed[1867],seed[1932],seed[4081],seed[2171],seed[3699],seed[3818],seed[3274],seed[2796],seed[1224],seed[172],seed[1267],seed[2641],seed[3646],seed[1893],seed[2990],seed[1262],seed[2943],seed[109],seed[1785],seed[2237],seed[2188],seed[108],seed[3942],seed[3775],seed[1740],seed[3859],seed[1051],seed[1292],seed[1567],seed[1031],seed[1836],seed[772],seed[3050],seed[1916],seed[2588],seed[2570],seed[1123],seed[3018],seed[1045],seed[287],seed[787],seed[1890],seed[1403],seed[3258],seed[1434],seed[931],seed[3284],seed[2715],seed[2994],seed[200],seed[3541],seed[2538],seed[1430],seed[72],seed[2565],seed[2844],seed[4038],seed[2885],seed[1165],seed[2836],seed[502],seed[59],seed[2154],seed[361],seed[1674],seed[3195],seed[1874],seed[20],seed[2215],seed[1772],seed[744],seed[869],seed[3507],seed[3974],seed[1088],seed[775],seed[3265],seed[1256],seed[2648],seed[1543],seed[188],seed[3918],seed[1767],seed[3402],seed[4077],seed[496],seed[3728],seed[1553],seed[1221],seed[490],seed[1842],seed[3148],seed[3551],seed[3980],seed[3320],seed[192],seed[3736],seed[2326],seed[3570],seed[2233],seed[2888],seed[3432],seed[1895],seed[2625],seed[2035],seed[1187],seed[3054],seed[3281],seed[1573],seed[3725],seed[2332],seed[444],seed[415],seed[688],seed[3594],seed[390],seed[2757],seed[413],seed[3826],seed[1317],seed[3075],seed[3709],seed[2606],seed[2179],seed[425],seed[2980],seed[3481],seed[2157],seed[3294],seed[1941],seed[345],seed[561],seed[1280],seed[892],seed[3058],seed[2117],seed[1053],seed[3987],seed[1186],seed[247],seed[2829],seed[2624],seed[1297],seed[48],seed[166],seed[2282],seed[1075],seed[1512],seed[3163],seed[955],seed[1451],seed[3383],seed[1231],seed[2449],seed[193],seed[312],seed[1036],seed[3595],seed[1961],seed[895],seed[473],seed[3738],seed[2724],seed[3630],seed[1499],seed[3863],seed[2969],seed[248],seed[3740],seed[2945],seed[1278],seed[2557],seed[1046],seed[875],seed[465],seed[2577],seed[1303],seed[249],seed[3791],seed[1617],seed[3864],seed[592],seed[3639],seed[3811],seed[451],seed[3463],seed[3529],seed[3187],seed[3620],seed[1597],seed[2192],seed[827],seed[1305],seed[659],seed[3223],seed[2044],seed[328],seed[3868],seed[3426],seed[3221],seed[958],seed[886],seed[436],seed[2181],seed[3210],seed[3707],seed[804],seed[1949],seed[1454],seed[2055],seed[388],seed[927],seed[252],seed[3785],seed[1701],seed[1537],seed[2516],seed[3549],seed[2629],seed[1655],seed[2095],seed[3522],seed[801],seed[3884],seed[1012],seed[684],seed[537],seed[3622],seed[3917],seed[770],seed[3453],seed[1098],seed[969],seed[3770],seed[3502],seed[3466],seed[2592],seed[2909],seed[3697],seed[693],seed[3504],seed[3889],seed[315],seed[1505],seed[3632],seed[633],seed[2195],seed[2890],seed[3136],seed[3002],seed[1448],seed[515],seed[1875],seed[1360],seed[3082],seed[3514],seed[2445],seed[1866],seed[3810],seed[3312],seed[2018],seed[2333],seed[1832],seed[3609],seed[3354],seed[1605],seed[3640],seed[1631],seed[2825],seed[210],seed[2750],seed[2300],seed[1275],seed[4086],seed[2223],seed[1557],seed[2307],seed[1983],seed[3053],seed[2948],seed[4095],seed[2512],seed[3298],seed[2291],seed[1862],seed[196],seed[1928],seed[867],seed[3324],seed[3220],seed[1716],seed[842],seed[3682],seed[2861],seed[877],seed[133],seed[482],seed[3579],seed[3706],seed[2628],seed[3370],seed[2871],seed[1523],seed[578],seed[3841],seed[2760],seed[3660],seed[1873],seed[769],seed[850],seed[4043],seed[1804],seed[2446],seed[2415],seed[3156],seed[1054],seed[1376],seed[3175],seed[703],seed[802],seed[2371],seed[765],seed[73],seed[3756],seed[69],seed[1489],seed[3858],seed[2367],seed[782],seed[321],seed[3914],seed[3144],seed[2499],seed[385],seed[2615],seed[1180],seed[2776],seed[2995],seed[3479],seed[2418],seed[2510],seed[1864],seed[2865],seed[3201],seed[1955],seed[3211],seed[1049],seed[1651],seed[3512],seed[585],seed[826],seed[1287],seed[2976],seed[640],seed[2848],seed[3543],seed[3036],seed[1978],seed[276],seed[1675],seed[517],seed[2152],seed[593],seed[851],seed[3157],seed[3247],seed[1626],seed[71],seed[2145],seed[768],seed[2459],seed[2014],seed[357],seed[1791],seed[2781],seed[3305],seed[897],seed[3028],seed[2312],seed[3411],seed[796],seed[3188],seed[3866],seed[1001],seed[1673],seed[156],seed[551],seed[3131],seed[3729],seed[2485],seed[1506],seed[2940],seed[3880],seed[2461],seed[300],seed[3951],seed[1632],seed[2753],seed[1940],seed[833],seed[1177],seed[1750],seed[3975],seed[191],seed[3510],seed[1338],seed[1869],seed[1061],seed[1527],seed[2121],seed[2193],seed[1421],seed[2169],seed[3382],seed[2711],seed[2401],seed[3717],seed[2464],seed[2110],seed[686],seed[2610],seed[574],seed[1758],seed[1226],seed[3705],seed[2944],seed[1733],seed[4027],seed[3259],seed[3118],seed[3442],seed[2794],seed[2103],seed[3996],seed[1811],seed[3523],seed[1880],seed[1126],seed[2092],seed[1713],seed[1406],seed[3552],seed[1229],seed[3553],seed[2281],seed[3056],seed[3485],seed[2733],seed[589],seed[2216],seed[3032],seed[2973],seed[3908],seed[813],seed[2346],seed[4045],seed[608],seed[3343],seed[1903],seed[745],seed[1560],seed[2151],seed[2907],seed[1821],seed[3369],seed[3425],seed[2642],seed[3856],seed[2806],seed[1566],seed[3012],seed[3840],seed[131],seed[3278],seed[1070],seed[513],seed[165],seed[1554],seed[1337],seed[1111],seed[268],seed[3698],seed[3431],seed[2132],seed[906],seed[1858],seed[122],seed[752],seed[634],seed[1485],seed[1948],seed[362],seed[476],seed[725],seed[2294],seed[2226],seed[1535],seed[1169],seed[1629],seed[2264],seed[2997],seed[1372],seed[3437],seed[3069],seed[0],seed[1906],seed[3048],seed[1004],seed[130],seed[177],seed[2868],seed[2849],seed[455],seed[1603],seed[577],seed[3174],seed[872],seed[3461],seed[3757],seed[1160],seed[23],seed[3506],seed[3153],seed[1008],seed[222],seed[2562],seed[1288],seed[937],seed[3132],seed[1578],seed[1339],seed[1072],seed[1795],seed[2703],seed[1319],seed[785],seed[1002],seed[3931],seed[3129],seed[1043],seed[1622],seed[3967],seed[2644],seed[4015],seed[4084],seed[125],seed[497],seed[1402],seed[2575],seed[1551],seed[2277],seed[1802],seed[3773],seed[3907],seed[4072],seed[1196],seed[761],seed[2342],seed[63],seed[3860],seed[3081],seed[1151],seed[2447],seed[1516],seed[2093],seed[571],seed[3396],seed[240],seed[259],seed[1924],seed[211],seed[2058],seed[3073],seed[3519],seed[4013],seed[1014],seed[3176],seed[2136],seed[136],seed[1175],seed[1323],seed[3779],seed[127],seed[2454],seed[1315],seed[2534],seed[3687],seed[3517],seed[2859],seed[2306],seed[2941],seed[3703],seed[555],seed[3766],seed[1184],seed[3219],seed[47],seed[2398],seed[1133],seed[3165],seed[2673],seed[3031],seed[184],seed[3629],seed[1140],seed[2419],seed[3286],seed[3711],seed[3801],seed[3429],seed[904],seed[4011],seed[2942],seed[3611],seed[4051],seed[2078],seed[2420],seed[460],seed[2573],seed[331],seed[3684],seed[3405],seed[1558],seed[1055],seed[1582],seed[3322],seed[2259],seed[1393],seed[1742],seed[2334],seed[2988],seed[1741],seed[563],seed[146],seed[212],seed[1593],seed[2275],seed[2187],seed[2545],seed[2252],seed[1640],seed[492],seed[1234],seed[378],seed[1418],seed[1702],seed[54],seed[982],seed[1780],seed[420],seed[1429],seed[3695],seed[3193],seed[560],seed[2402],seed[433],seed[2579],seed[4006],seed[631],seed[1074],seed[458],seed[3566],seed[2348],seed[1225],seed[1926],seed[1824],seed[2175],seed[2205],seed[3057],seed[876],seed[475],seed[2939],seed[3591],seed[1747],seed[1479],seed[1199],seed[1057],seed[3470],seed[2820],seed[2896],seed[2357],seed[2809],seed[3748],seed[2714],seed[3403],seed[2126],seed[2470],seed[1953],seed[2857],seed[901],seed[152],seed[3052],seed[4063],seed[3114],seed[1820],seed[3804],seed[2427],seed[2572],seed[4076],seed[1810],seed[1946],seed[2482],seed[3072],seed[1086],seed[1266],seed[1179],seed[1845],seed[479],seed[1913],seed[1085],seed[3349],seed[3955],seed[2837],seed[864],seed[2792],seed[3491],seed[705],seed[3406],seed[422],seed[3776],seed[3751],seed[456],seed[1296],seed[2555],seed[1781],seed[30],seed[3539],seed[1760],seed[2397],seed[15],seed[3790],seed[650],seed[2109],seed[929],seed[2766],seed[3143],seed[844],seed[3842],seed[2020],seed[941],seed[548],seed[3525],seed[2383],seed[911],seed[2782],seed[2901],seed[648],seed[2893],seed[620],seed[3598],seed[2543],seed[2303],seed[3896],seed[737],seed[3364],seed[3366],seed[2238],seed[1093],seed[25],seed[3159],seed[2255],seed[2327],seed[3575],seed[2159],seed[2762],seed[999],seed[3799],seed[1309],seed[1089],seed[697],seed[2356],seed[535],seed[3422],seed[528],seed[3380],seed[1990],seed[2951],seed[2731],seed[2950],seed[2877],seed[846],seed[2826],seed[843],seed[2904],seed[3750],seed[572],seed[147],seed[3822],seed[3845],seed[1515],seed[1530],seed[1524],seed[1040],seed[794],seed[2403],seed[3218],seed[3661],seed[2304],seed[3784],seed[2827],seed[3040],seed[151],seed[3151],seed[598],seed[1128],seed[748],seed[933],seed[3152],seed[499],seed[1801],seed[670],seed[3068],seed[2011],seed[776],seed[3496],seed[1730],seed[2897],seed[2274],seed[2571],seed[557],seed[1340],seed[1343],seed[2779],seed[296],seed[3623],seed[1320],seed[195],seed[3145],seed[2991],seed[3716],seed[3280],seed[3059],seed[1080],seed[2536],seed[2494],seed[730],seed[2513],seed[223],seed[443],seed[132],seed[1991],seed[2883],seed[3020],seed[1495],seed[3226],seed[1989],seed[3981],seed[1058],seed[3733],seed[2165],seed[2899],seed[3587],seed[1829],seed[4031],seed[2996],seed[584],seed[1789],seed[2056],seed[3460],seed[1498],seed[2341],seed[2040],seed[273],seed[1703],seed[3293],seed[2667],seed[625],seed[2884],seed[2852],seed[3999],seed[3540],seed[2585],seed[2359],seed[1644],seed[2484],seed[797],seed[1130],seed[2474],seed[2460],seed[3771],seed[3596],seed[3528],seed[1678],seed[3438],seed[194],seed[3638],seed[186],seed[1541],seed[565],seed[2881],seed[617],seed[531],seed[1386],seed[3829],seed[4046],seed[1082],seed[3351],seed[638],seed[820],seed[3870],seed[3046],seed[143],seed[1725],seed[372],seed[3589],seed[3936],seed[2959],seed[511],seed[1611],seed[414],seed[2353],seed[2646],seed[3416],seed[3106],seed[141],seed[4080],seed[540],seed[3212],seed[2926],seed[526],seed[1380],seed[2501],seed[3887],seed[3352],seed[3902],seed[438],seed[175],seed[2290],seed[3869],seed[1475],seed[3026],seed[809],seed[2207],seed[3608],seed[1428],seed[1956],seed[1302],seed[66],seed[189],seed[3749],seed[2451],seed[3030],seed[307],seed[2128],seed[2072],seed[2329],seed[4036],seed[2804],seed[712],seed[951],seed[3166],seed[1779],seed[3169],seed[3546],seed[1788],seed[1193],seed[3098],seed[812],seed[167],seed[2086],seed[233],seed[2479],seed[4055],seed[3696],seed[2748],seed[3332],seed[472],seed[1211],seed[4003],seed[3229],seed[1414],seed[2561],seed[2472],seed[3445],seed[2962],seed[3806],seed[1634],seed[583],seed[3242],seed[2288],seed[1571],seed[3585],seed[3358],seed[848],seed[3605],seed[524],seed[3946],seed[665],seed[3774],seed[2594],seed[3389],seed[256],seed[343],seed[509],seed[1382],seed[1529],seed[2065],seed[2395],seed[2957],seed[1777],seed[3164],seed[1695],seed[1840],seed[1148],seed[3409],seed[2085],seed[3817],seed[351],seed[1107],seed[3267],seed[788],seed[790],seed[815],seed[2314],seed[2296],seed[2631],seed[1507],seed[3126],seed[3296],seed[2887],seed[742],seed[503],seed[898],seed[3302],seed[3904],seed[60],seed[754],seed[859],seed[3300],seed[3788],seed[139],seed[1528],seed[2468],seed[3557],seed[1400],seed[1459],seed[1723],seed[3340],seed[1959],seed[1350],seed[689],seed[2704],seed[2919],seed[1387],seed[3927],seed[2999],seed[3890],seed[2993],seed[2863],seed[402],seed[3943],seed[1015],seed[2316],seed[1104],seed[169],seed[1252],seed[1714],seed[2146],seed[1011],seed[2050],seed[520],seed[3319],seed[3653],seed[2203],seed[3824],seed[408],seed[1440],seed[2791],seed[145],seed[1009],seed[1671],seed[2089],seed[106],seed[1531],seed[1006],seed[4016],seed[236],seed[1446],seed[3237],seed[2037],seed[784],seed[675],seed[914],seed[1910],seed[1969],seed[1784],seed[3787],seed[3702],seed[3093],seed[450],seed[3724],seed[3601],seed[439],seed[1927],seed[971],seed[542],seed[915],seed[1915],seed[10],seed[1154],seed[1646],seed[1743],seed[3882],seed[1463],seed[17],seed[1132],seed[943],seed[176],seed[916],seed[2564],seed[1584],seed[1883],seed[395],seed[3084],seed[3586],seed[1766],seed[1871],seed[2478],seed[107],seed[1149],seed[2133],seed[266],seed[564],seed[3550],seed[3667],seed[1171],seed[3920],seed[2839],seed[3230],seed[1720],seed[454],seed[3337],seed[2535],seed[1341],seed[1468],seed[2183],seed[2311],seed[1805],seed[3582],seed[1793],seed[1114],seed[599],seed[2438],seed[957],seed[310],seed[392],seed[3686],seed[1771],seed[3374],seed[1888],seed[3109],seed[749],seed[1493],seed[4079],seed[4017],seed[1947],seed[1162],seed[4029],seed[701],seed[82],seed[4020],seed[3011],seed[2135],seed[3997],seed[1250],seed[3618],seed[1583],seed[1694],seed[3808],seed[3819],seed[2866],seed[913],seed[397],seed[657],seed[3231],seed[821],seed[3743],seed[1467],seed[1904],seed[3958],seed[374],seed[4040],seed[3655],seed[1565],seed[3592],seed[3534],seed[3578],seed[2666],seed[2176],seed[1469],seed[3034],seed[421],seed[1259],seed[2396],seed[1778],seed[1884],seed[3669],seed[1163],seed[2394],seed[3657],seed[1677],seed[695],seed[126],seed[2261],seed[2604],seed[739],seed[1425],seed[3149],seed[2688],seed[2713],seed[2015],seed[118],seed[1988],seed[1419],seed[1828],seed[2210],seed[2652],seed[1084],seed[2355],seed[549],seed[1146],seed[2789],seed[2636],seed[740],seed[2201],seed[65],seed[1581],seed[350],seed[1216],seed[2645],seed[1851],seed[924],seed[2305],seed[2217],seed[3966],seed[4064],seed[3827],seed[1660],seed[3088],seed[2410],seed[3972],seed[1841],seed[1735],seed[587],seed[4085],seed[1473],seed[3180],seed[921],seed[2786],seed[28],seed[871],seed[1717],seed[2041],seed[3234],seed[2721],seed[434],seed[3111],seed[3041],seed[639],seed[2684],seed[3039],seed[3580],seed[1876],seed[2345],seed[644],seed[3117],seed[3531],seed[2405],seed[1023],seed[3001],seed[905],seed[3617],seed[387],seed[2254],seed[2424],seed[4073],seed[3225],seed[1487],seed[1757],seed[405],seed[3303],seed[3271],seed[3713],seed[37],seed[1397],seed[3588],seed[3726],seed[2569],seed[750],seed[1290],seed[3295],seed[2700],seed[807],seed[2680],seed[124],seed[3603],seed[1786],seed[1143],seed[359],seed[1105],seed[398],seed[340],seed[3719],seed[3100],seed[1318],seed[2349],seed[1257],seed[3912],seed[1938],seed[3915],seed[1245],seed[618],seed[2986],seed[76],seed[3547],seed[3228],seed[1905],seed[573],seed[2477],seed[3710],seed[3019],seed[681],seed[1092],seed[2491],seed[404],seed[3763],seed[1511],seed[228],seed[171],seed[727],seed[3542],seed[271],seed[677],seed[3025],seed[1638],seed[1359],seed[2368],seed[3318],seed[239],seed[746],seed[1488],seed[493],seed[3834],seed[3913],seed[708],seed[2799],seed[3768],seed[2036],seed[2229],seed[1304],seed[1534],seed[3634],seed[1598],seed[1768],seed[3988],seed[2400],seed[3621],seed[508],seed[3350],seed[2921],seed[384],seed[3077],seed[3664],seed[2755],seed[1798],seed[2105],seed[3903],seed[498],seed[658],seed[44],seed[3015],seed[3922],seed[373],seed[635],seed[1698],seed[2741],seed[1547],seed[1328],seed[1020],seed[2235],seed[1144],seed[3139],seed[2267],seed[1732],seed[324],seed[1753],seed[830],seed[1150],seed[3497],seed[39],seed[1066],seed[309],seed[2956],seed[3637],seed[487],seed[170],seed[3244],seed[3083],seed[3137],seed[3215],seed[1147],seed[481],seed[1982],seed[566],seed[2747],seed[3894],seed[2580],seed[3116],seed[1687],seed[2966],seed[2635],seed[2313],seed[1330],seed[2623],seed[462],seed[882],seed[217],seed[3720],seed[320],seed[2481],seed[1235],seed[968],seed[3256],seed[3119],seed[3830],seed[393],seed[3270],seed[731],seed[1447],seed[3888],seed[43],seed[758],seed[974],seed[2930],seed[2683],seed[483],seed[629],seed[988],seed[2240],seed[1490],seed[2891],seed[2278],seed[2697],seed[2366],seed[3835],seed[3919],seed[3604],seed[2874],seed[3217],seed[2931],seed[255],seed[2158],seed[2271],seed[806],seed[52],seed[994],seed[250],seed[1650],seed[1613],seed[3607],seed[1415],seed[1413],seed[1206],seed[2178],seed[683],seed[500],seed[3521],seed[506],seed[291],seed[3167],seed[1321],seed[2875],seed[45],seed[2964],seed[1356],seed[3078],seed[3984],seed[1029],seed[1596],seed[2450],seed[3559],seed[1748],seed[2337],seed[2272],seed[2797],seed[2344],seed[2596],seed[2695],seed[158],seed[4053],seed[1708],seed[2012],seed[3873],seed[2710],seed[2352],seed[2031],seed[2719],seed[926],seed[1228],seed[559],seed[491],seed[2894],seed[1846],seed[3619],seed[803],seed[2429],seed[1033],seed[1332],seed[3932],seed[2489],seed[1135],seed[3346],seed[2612],seed[2522],seed[2739],seed[1974],seed[1594],seed[3197],seed[3173],seed[2389],seed[1354],seed[1039],seed[856],seed[2033],seed[1960],seed[2862],seed[721],seed[3769],seed[3558],seed[2622],seed[902],seed[919],seed[3357],seed[2589],seed[153],seed[3367],seed[651],seed[3456],seed[3606],seed[959],seed[2856],seed[3459],seed[1542],seed[49],seed[4047],seed[3395],seed[4035],seed[85],seed[278],seed[1478],seed[3755],seed[168],seed[2375],seed[148],seed[369],seed[1426],seed[614],seed[245],seed[3962],seed[1633],seed[488],seed[4],seed[2581],seed[837],seed[2679],seed[2098],seed[1822],seed[347],seed[2005],seed[610],seed[3708],seed[3133],seed[981],seed[103],seed[2758],seed[1630],seed[2431],seed[3398],seed[1661],seed[3199],seed[308],seed[1286],seed[1901],seed[2851],seed[1664],seed[698],seed[1207],seed[3042],seed[2526],seed[46],seed[1849],seed[117],seed[2685],seed[1881],seed[2250],seed[3440],seed[1116],seed[3063],seed[3956],seed[1679],seed[1657],seed[3959],seed[2437],seed[1272],seed[868],seed[3208],seed[2847],seed[3421],seed[2915],seed[755],seed[2066],seed[1432],seed[2725],seed[2798],seed[218],seed[2189],seed[3467],seed[83],seed[3691],seed[3615],seed[1996],seed[3372],seed[4052],seed[2870],seed[3681],seed[3625],seed[910],seed[522],seed[3064],seed[2832],seed[1522],seed[87],seed[558],seed[702],seed[655],seed[2488],seed[411],seed[977],seed[98],seed[3986],seed[896],seed[2582],seed[474],seed[3765],seed[2780],seed[9],seed[2503],seed[3926],seed[1686],seed[162],seed[2992],seed[3251],seed[3209],seed[586],seed[2],seed[3690],seed[2273],seed[2933],seed[2961],seed[1830],seed[2074],seed[4082],seed[2726],seed[437],seed[1101],seed[976],seed[12],seed[99],seed[1158],seed[3561],seed[2563],seed[1609],seed[764],seed[105],seed[847],seed[226],seed[1295],seed[3263],seed[1247],seed[401],seed[1112],seed[964],seed[3368],seed[2480],seed[3745],seed[1159],seed[1680],seed[3954],seed[67],seed[2360],seed[2323],seed[34],seed[2161],seed[3780],seed[2293],seed[1999],seed[3150],seed[3115],seed[3742],seed[2234],seed[1872],seed[2508],seed[3654],seed[3384],seed[417],seed[406],seed[3317],seed[4050],seed[1188],seed[2407],seed[1125],seed[607],seed[2506],seed[2096],seed[950],seed[831],seed[197],seed[3732],seed[2559],seed[2978],seed[962],seed[2821],seed[3635],seed[3851],seed[2675],seed[3359],seed[3375],seed[2817],seed[79],seed[2546],seed[1591],seed[280],seed[3158],seed[2131],seed[2614],seed[2527],seed[2317],seed[1007],seed[3449],seed[2947],seed[1763],seed[2197],seed[2309],seed[3929],seed[1361],seed[747],seed[2689],seed[2960],seed[3569],seed[3016],seed[1917],seed[1852],seed[612],seed[1800],seed[711],seed[461],seed[2900],seed[383],seed[137],seed[2184],seed[2463],seed[1833],seed[1333],seed[282],seed[760],seed[3476],seed[292],seed[1357],seed[2227],seed[3644],seed[2245],seed[2315],seed[3567],seed[900],seed[3891],seed[346],seed[1976],seed[1658],seed[3797],seed[41],seed[3257],seed[3701],seed[1255],seed[1076],seed[909],seed[2139],seed[1138],seed[580],seed[1311],seed[3815],seed[3998],seed[2452],seed[1018],seed[2059],seed[1243],seed[2946],seed[1377],seed[3941],seed[1608],seed[284],seed[3793],seed[2285],seed[2208],seed[1620],seed[2114],seed[539],seed[2983],seed[2749],seed[2283],seed[3648],seed[2289],seed[925],seed[1050],seed[1293],seed[1751],seed[3683],seed[3680],seed[4004],seed[2640],seed[1482],seed[1131],seed[3849],seed[3626],seed[3233],seed[3009],seed[3189],seed[3833],seed[237],seed[116],seed[33],seed[51],seed[2542],seed[3995],seed[1503],seed[2770],seed[3005],seed[3792],seed[4008],seed[1826],seed[1886],seed[4058],seed[2340],seed[2910],seed[1019],seed[2232],seed[92],seed[330],seed[3939],seed[2935],seed[2765],seed[2505],seed[1971],seed[2660],seed[3862],seed[3832],seed[2761],seed[653],seed[3253],seed[3933],seed[3102],seed[1726],seed[341],seed[1355],seed[979],seed[2358],seed[1263],seed[619],seed[3194],seed[1706],seed[1083],seed[432],seed[1992],seed[2191],seed[2043],seed[2708],seed[2558],seed[1770],seed[453],seed[1178],seed[2544],seed[2123],seed[1450],seed[2118],seed[1232],seed[2045],seed[2231],seed[2213],seed[3854],seed[2917],seed[570],seed[21],seed[1683],seed[3688],seed[3183],seed[1065],seed[3435],seed[3415],seed[836],seed[1589],seed[2286],seed[3934],seed[1063],seed[3490],seed[3970],seed[1041],seed[814],seed[829],seed[3642],seed[932],seed[810],seed[1625],seed[792],seed[1607],seed[3004],seed[1891],seed[2672],seed[2302],seed[756],seed[1755],seed[2029],seed[3043],seed[2369],seed[736],seed[4056],seed[1604],seed[2433],seed[1847],seed[2705],seed[2734],seed[270],seed[3092],seed[2912],seed[283],seed[3612],seed[1856],seed[2476],seed[2858],seed[2785],seed[3283],seed[2663],seed[2905],seed[1616],seed[2590],seed[3455],seed[2702],seed[3419],seed[2025],seed[884],seed[3472],seed[1574],seed[1642],seed[533],seed[2754],seed[3014],seed[2764],seed[543],seed[2225],seed[728],seed[2583],seed[879],seed[2101],seed[1021],seed[1168],seed[918],seed[3649],seed[538],seed[1564],seed[1056],seed[1759],seed[1705],seed[4092],seed[1456],seed[3568],seed[2143],seed[3205],seed[2462],seed[2243],seed[2613],seed[2370],seed[707],seed[2443],seed[1170],seed[1980],seed[779],seed[135],seed[2063],seed[1544],seed[187],seed[3241],seed[3436],seed[2046],seed[2952],seed[3679],seed[3177],seed[2658],seed[262],seed[1003],seed[1268],seed[1152],seed[2330],seed[2639],seed[2198],seed[2413],seed[1662],seed[1472],seed[1395],seed[164],seed[1807],seed[823],seed[2846],seed[3309],seed[96],seed[2321],seed[723],seed[673],seed[2090],seed[716],seed[656],seed[2144],seed[2694],seed[1769],seed[2112],seed[1283],seed[1237],seed[3731],seed[2554],seed[3982],seed[2385],seed[1920],seed[832],seed[1525],seed[956],seed[636],seed[4091],seed[285],seed[3447],seed[1555],seed[1970],seed[1639],seed[936],seed[2822],seed[1823],seed[1265],seed[609],seed[1827],seed[1692],seed[3345],seed[2172],seed[337],seed[3272],seed[1615],seed[1612],seed[3508],seed[3899],seed[2584],seed[2038],seed[883],seed[3338],seed[1722],seed[3573],seed[996],seed[3138],seed[1587],seed[322],seed[3101],seed[972],seed[2932],seed[3124],seed[1127],seed[91],seed[1017],seed[726],seed[3944],seed[459],seed[2953],seed[628],seed[1814],seed[2740],seed[2001],seed[3344],seed[2148],seed[2654],seed[3067],seed[281],seed[2265],seed[2752],seed[778],seed[3090],seed[2855],seed[2416],seed[3636],seed[1684],seed[863],seed[269],seed[1307],seed[3965],seed[3390],seed[3747],seed[3323],seed[2391],seed[3376],seed[1973],seed[198],seed[2840],seed[3045],seed[2280],seed[3182],seed[2968],seed[2763],seed[983],seed[1649],seed[2019],seed[265],seed[3548],seed[1059],seed[1669],seed[3712],seed[1067],seed[3831],seed[1838],seed[2399],seed[2609],seed[3692],seed[2818],seed[3154],seed[1517],seed[2669],seed[354],seed[3689],seed[3356],seed[389],seed[1399],seed[1457],seed[1572],seed[2387],seed[3037],seed[1621],seed[2174],seed[2498],seed[2963],seed[2872],seed[2574],seed[3495],seed[1433],seed[3898],seed[1546],seed[2934],seed[2469],seed[2032],seed[1809],seed[2196],seed[992],seed[3600],seed[514],seed[714],seed[183],seed[2325],seed[3107],seed[3140],seed[3450],seed[111],seed[771],seed[920],seed[1254],seed[2743],seed[3289],seed[970],seed[3299],seed[3990],seed[2618],seed[3171],seed[3878],seed[3532],seed[2129],seed[1052],seed[3439],seed[1889],seed[889],seed[504],seed[2119],seed[364],seed[1367],seed[306],seed[3584],seed[3204],seed[4054],seed[822],seed[370],seed[3314],seed[1212],seed[2435],seed[2751],seed[3168],seed[2716],seed[1729],seed[1986],seed[2729],seed[3315],seed[3412],seed[261],seed[3857],seed[1069],seed[4078],seed[547],seed[3816],seed[1198],seed[2655],seed[3994],seed[3960],seed[1995],seed[2047],seed[1958],seed[295],seed[4012],seed[3091],seed[3400],seed[1000],seed[264],seed[1427],seed[1124],seed[562],seed[3501],seed[594],seed[1203],seed[1253],seed[2116],seed[2637],seed[154],seed[980],seed[2257],seed[1412],seed[3482],seed[3473],seed[732],seed[3694],seed[2153],seed[1627],seed[2674],seed[1269],seed[2351],seed[1389],seed[2166],seed[1392],seed[3576],seed[2981],seed[4039],seed[352],seed[2262],seed[3477],seed[26],seed[2511],seed[1962],seed[3062],seed[316],seed[3825],seed[2336],seed[1274],seed[1641],seed[1194],seed[215],seed[2379],seed[2647],seed[3393],seed[3408],seed[144],seed[3511],seed[2287],seed[1563],seed[928],seed[3122],seed[1273],seed[3307],seed[62],seed[3500],seed[201],seed[1911],seed[2319],seed[2732],seed[2718],seed[1939],seed[1081],seed[2914],seed[1480],seed[3821],seed[214],seed[1853],seed[3335],seed[2744],seed[1022],seed[2458],seed[1994],seed[3292],seed[3783],seed[3807],seed[2717],seed[4088],seed[104],seed[3488],seed[3693],seed[912],seed[2682],seed[4000],seed[263],seed[1032],seed[1176],seed[2595],seed[874],seed[3021],seed[2414],seed[1984],seed[780],seed[2099],seed[632],seed[138],seed[3761],seed[3530],seed[2568],seed[569],seed[2841],seed[1998],seed[3852],seed[2879],seed[3287],seed[1455],seed[1737],seed[3746],seed[3897],seed[2266],seed[2211],seed[14],seed[1102],seed[334],seed[2268],seed[1783],seed[507],seed[2607],seed[3252],seed[3803],seed[1854],seed[363],seed[2392],seed[3647],seed[1383],seed[2845],seed[1817],seed[3076],seed[379],seed[2529],seed[478],seed[1552],seed[19],seed[3916],seed[1665],seed[1600],seed[1445],seed[1349],seed[1700],seed[2814],seed[2989],seed[1486],seed[3007],seed[3110],seed[965],seed[2892],seed[323],seed[3254],seed[1937],seed[800],seed[1504],seed[4014],seed[3103],seed[603],seed[1120],seed[907],seed[2880],seed[1197],seed[2256],seed[1610],seed[944],seed[2120],seed[179],seed[3483],seed[1028],seed[4032],seed[1727],seed[3554],seed[1746],seed[3938],seed[942],seed[1586],seed[234],seed[1559],seed[2500],seed[2578],seed[484],seed[2771],seed[3715],seed[3160],seed[1371],seed[3855],seed[3651],seed[3505],seed[3645],seed[1844],seed[2502],seed[1261],seed[2298],seed[530],seed[3373],seed[2269],seed[74],seed[333],seed[3250],seed[1954],seed[3678],seed[1799],seed[2067],seed[3658],seed[849],seed[2911],seed[1711],seed[3814],seed[3652],seed[394],seed[3261],seed[3973],seed[1270],seed[1164],seed[3992],seed[1182],seed[3097],seed[205],seed[2677],seed[2170],seed[3249],seed[140],seed[428],seed[3969],seed[3430],seed[1606],seed[110],seed[1064],seed[409],seed[3730],seed[2062],seed[2634],seed[2854],seed[947],seed[299],seed[114],seed[1520],seed[182],seed[2998],seed[3222],seed[2549],seed[246],seed[329],seed[3650],seed[3207],seed[3509],seed[2324],seed[1209],seed[2520],seed[1481],seed[2361],seed[275],seed[2057],seed[2013],seed[468],seed[1190],seed[1129],seed[1411],seed[1260],seed[568],seed[2530],seed[2111],seed[1294],seed[687],seed[469],seed[1957],seed[431],seed[2515],seed[1819],seed[691],seed[3232],seed[3964],seed[880],seed[2601],seed[178],seed[3434],seed[1908],seed[786],seed[2657],seed[805],seed[2068],seed[2617],seed[1218],seed[3820],seed[2805],seed[4026],seed[1460],seed[1204],seed[1435],seed[1024],seed[2728],seed[3413],seed[2916],seed[2204],seed[3392],seed[2838],seed[181],seed[2404],seed[1929],seed[2200],seed[1313],seed[3562],seed[1142],seed[1483],seed[423],seed[3924],seed[3443],seed[1690],seed[1035],seed[505],seed[2816],seed[2665],seed[774],seed[4049],seed[2735],seed[2547],seed[1569],seed[1443],seed[2382],seed[984],seed[1987],seed[88],seed[1244],seed[841],seed[987],seed[3759],seed[358],seed[1774],seed[1602],seed[525],seed[2597],seed[400],seed[4048],seed[2643],seed[3262],seed[704],seed[3752],seed[674],seed[2775],seed[1979],seed[1935],seed[2651],seed[3910],seed[3288],seed[2260],seed[3044],seed[516],seed[35],seed[2007],seed[150],seed[1985],seed[855],seed[3739],seed[862],seed[2670],seed[2457],seed[3850],seed[903],seed[1477],seed[3074],seed[789],seed[327],seed[2727],seed[1636],seed[3671],seed[311],seed[1369],seed[3672],seed[3662],seed[78],seed[2599],seed[3094],seed[873],seed[2556],seed[2737],seed[2552],seed[3753],seed[1496],seed[3457],seed[2707],seed[3125],seed[1754],seed[1298],seed[1351],seed[317],seed[466],seed[3027],seed[3087],seed[2378],seed[1097],seed[3949],seed[1739],seed[1335],seed[1526],seed[3876],seed[2698],seed[1401],seed[3404],seed[1205],seed[2514],seed[3564],seed[899],seed[480],seed[209],seed[4090],seed[1712],seed[3828],seed[678],seed[2955],seed[1718],seed[2690],seed[1704],seed[865],seed[1601],seed[2028],seed[3722],seed[2440],seed[1462],seed[3754],seed[2807],seed[3853],seed[3070],seed[2372],seed[767],seed[2709],seed[1812],seed[3794],seed[2426],seed[1217],seed[2276],seed[2860],seed[3475],seed[2678],seed[1775],seed[1342],seed[3035],seed[2850],seed[2490],seed[2745],seed[2363],seed[2475],seed[1436],seed[1652],seed[3581],seed[3361],seed[3095],seed[819],seed[3360],seed[2228],seed[2746],seed[1925],seed[3487],seed[303],seed[1590],seed[1691],seed[3844],seed[1707],seed[2455],seed[1635],seed[2813],seed[791],seed[180],seed[934],seed[1818],seed[2808],seed[2075],seed[2083],seed[272],seed[2155],seed[1037],seed[452],seed[2466],seed[289],seed[3555],seed[751],seed[2519],seed[294],seed[606],seed[3130],seed[3494],seed[2423],seed[2898],seed[709],seed[349],seed[2122],seed[120],seed[3484],seed[4093],seed[3146],seed[816],seed[3333],seed[3577],seed[2331],seed[2456],seed[1562],seed[3128],seed[3071],seed[1258],seed[738],seed[61],seed[649],seed[2308],seed[216],seed[1416],seed[4019],seed[923],seed[1157],seed[1899],seed[3885],seed[2149],seed[3216],seed[998],seed[3989],seed[3336],seed[3433],seed[319],seed[2027],seed[1264],seed[68],seed[1281],seed[672],seed[1685],seed[596],seed[799],seed[326],seed[1249],seed[3474],seed[161],seed[2975],seed[3310],seed[930],seed[2428],seed[3381],seed[940],seed[866],seed[510],seed[3524],seed[3414],seed[2493],seed[2800],seed[3134],seed[3823],seed[2611],seed[1967],seed[3945],seed[24],seed[2087],seed[2687],seed[954],seed[1016],seed[3423],seed[2365],seed[3000],seed[2742],seed[1936],seed[1997],seed[637],seed[1538],seed[3008],seed[3179],seed[2783],seed[3940],seed[1471],seed[3112],seed[1172],seed[1417],seed[1223],seed[2539],seed[3326],seed[3363],seed[3613],seed[604],seed[2364],seed[1628],seed[3947],seed[818],seed[613],seed[4028],seed[3796],seed[1444],seed[2377],seed[3113],seed[1381],seed[3266],seed[206],seed[1857],seed[783],seed[3033],seed[2186],seed[3424],seed[4062],seed[1238],seed[512],seed[1122],seed[5],seed[220],seed[1902],seed[1167],seed[2081],seed[84],seed[1894],seed[22],seed[494],seed[1756],seed[4001],seed[1113],seed[3468],seed[2060],seed[2134],seed[2249],seed[2000],seed[2284],seed[2824],seed[2140],seed[1378],seed[948],seed[3843],seed[1548],seed[3135],seed[1580],seed[1213],seed[1912],seed[1792],seed[251],seed[3198],seed[2064],seed[840],seed[2002],seed[2310],seed[1345],seed[845],seed[534],seed[2322],seed[2843],seed[2889],seed[1096],seed[995],seed[2603],seed[2194],seed[1161],seed[254],seed[298],seed[4030],seed[1697],seed[3486],seed[3089],seed[2819],seed[55],seed[377],seed[2496],seed[3781],seed[1236],seed[260],seed[1681],seed[890],seed[2938],seed[3418],seed[36],seed[32],seed[3304],seed[1539],seed[1568],seed[1241],seed[360],seed[2659],seed[1423],seed[2242],seed[1922],seed[743],seed[2936],seed[2039],seed[3493],seed[2082],seed[682],seed[3297],seed[1721],seed[757],seed[1592],seed[3921],seed[2388],seed[314],seed[3925],seed[2073],seed[290],seed[2518],seed[852],seed[2320],seed[3277],seed[3991],seed[227],seed[1532],seed[396],seed[258],seed[1859],seed[2965],seed[949],seed[2925],seed[1951],seed[2292],seed[1422],seed[2949],seed[3627],seed[366],seed[1476],seed[447],seed[1710],seed[1863],seed[601],seed[661],seed[3099],seed[1347],seed[1300],seed[1322],seed[3778],seed[2010],seed[3017],seed[1808],seed[835],seed[1848],seed[627],seed[1312],seed[1659],seed[2248],seed[667],seed[3536],seed[1667],seed[27],seed[2873],seed[2104],seed[766],seed[2448],seed[654],seed[2219],seed[2830],seed[355],seed[1752],seed[448],seed[2160],seed[365],seed[3196],seed[1325],seed[706],seed[3331],seed[427],seed[3362],seed[1156],seed[1110],seed[1868],seed[3162],seed[2202],seed[3704],seed[121],seed[1963],seed[2650],seed[1437],seed[3471],seed[3616],seed[4057],seed[2053],seed[1474],seed[3723],seed[1595],seed[3928],seed[399],seed[2630],seed[3085],seed[2142],seed[1787],seed[3838],seed[3282],seed[722],seed[878],seed[1222],seed[3677],seed[1484],seed[3812],seed[149],seed[3224],seed[1764],seed[1508],seed[2220],seed[2301],seed[616],seed[204],seed[119],seed[2693],seed[1839],seed[1470],seed[1410],seed[2902],seed[2354],seed[734],seed[1897],seed[1215],seed[735],seed[3161],seed[230],seed[3328],seed[2720],seed[666],seed[860],seed[2886],seed[1513],seed[3560],seed[2077],seed[2214],seed[185],seed[985],seed[58],seed[3239],seed[305],seed[3410],seed[1825],seed[3777],seed[1981],seed[3308],seed[1174],seed[1358],seed[3458],seed[3245],seed[1242],seed[546],seed[2773],seed[3685],seed[2106],seed[3673],seed[477],seed[2137],seed[446],seed[1137],seed[1119],seed[3633],seed[3985],seed[416],seed[2026],seed[163],seed[893],seed[3979],seed[2927],seed[2224],seed[3371],seed[2156],seed[1299],seed[412],seed[208],seed[102],seed[2533],seed[2924],seed[1952],seed[3758],seed[2124],seed[3744],seed[1588],seed[1],seed[336],seed[2869],seed[3255],seed[2439],seed[2828],seed[1336],seed[221],seed[3656],seed[3061],seed[495],seed[2523],seed[1087],seed[3837],seed[1918],seed[2633],seed[224],seed[1219],seed[2795],seed[3451],seed[2417],seed[692],seed[2920],seed[3334],seed[3798],seed[1166],seed[3023],seed[660],seed[602],seed[1060],seed[811],seed[1944],seed[1579],seed[1452],seed[2147],seed[2509],seed[527],seed[2328],seed[4005],seed[1277],seed[643],seed[1071],seed[2668],seed[332],seed[2738],seed[2069],seed[1090],seed[3185],seed[257],seed[1797],seed[1734],seed[1696],seed[1914],seed[1656],seed[2586],seed[1407],seed[645],seed[1115],seed[1047],seed[2246],seed[1724],seed[1103],seed[2023],seed[3060],seed[579],seed[1136],seed[2138],seed[2006],seed[1536],seed[908],seed[2239],seed[1062],seed[3968],seed[4024],seed[2408],seed[94],seed[857],seed[541],seed[588],seed[2541],seed[441],seed[3327],seed[710],seed[2335],seed[1306],seed[3923],seed[1898],seed[86],seed[3846],seed[2182],seed[2548],seed[1834],seed[1108],seed[442],seed[418],seed[1314],seed[2768],seed[501],seed[2835],seed[1271],seed[2810],seed[3273],seed[2793],seed[3883],seed[664],seed[2190],seed[3847],seed[356],seed[1749],seed[241],seed[2985],seed[1034],seed[2723],seed[2163],seed[3142],seed[824],seed[939],seed[2895],seed[2421],seed[3489],seed[1042],seed[3243],seed[277],seed[3190],seed[1934],seed[2049],seed[3051],seed[3670],seed[3013],seed[3556],seed[825],seed[798],seed[1200],seed[2071],seed[3565],seed[715],seed[2903],seed[891],seed[4007],seed[1835],seed[242],seed[338],seed[3503],seed[3737],seed[93],seed[1738],seed[4089],seed[1500],seed[621],seed[1492],seed[3417],seed[2409],seed[1373],seed[2712],seed[2487],seed[1648],seed[267],seed[1663],seed[3246],seed[1645],seed[2374],seed[1765],seed[935],seed[2164],seed[4069],seed[3772],seed[3735],seed[403],seed[225],seed[1877],seed[4023],seed[13],seed[1892],seed[3782],seed[3105],seed[3545],seed[3341],seed[4068],seed[1831],seed[2878],seed[3452],seed[3120],seed[1118],seed[1348],seed[1326],seed[2971],seed[2467],seed[3533],seed[1449],seed[81],seed[615],seed[3498],seed[1285],seed[391],seed[3665],seed[3276],seed[3516],seed[2802],seed[3170],seed[279],seed[741],seed[3428],seed[2177],seed[1282],seed[3909],seed[3055],seed[440],seed[817],seed[1668],seed[1431],seed[2212],seed[4044],seed[293],seed[3886],seed[556],seed[1424],seed[3628],seed[2411],seed[2373],seed[4071],seed[2030],seed[1374],seed[1331],seed[2567],seed[232],seed[3200],seed[986],seed[2209],seed[57],seed[626],seed[3394],seed[519],seed[2434],seed[2620],seed[1943],seed[449],seed[759],seed[2042],seed[2598],seed[157],seed[630],seed[1715],seed[3911],seed[1699],seed[174],seed[1141],seed[1079],seed[3446],seed[1619],seed[3108],seed[2384],seed[75],seed[2094],seed[70],seed[2778],seed[1191],seed[978],seed[3227],seed[2270],seed[2815],seed[3900],seed[1790],seed[2222],seed[2662],seed[3248],seed[3721],seed[4042],seed[3397],seed[2653],seed[3339],seed[3593],seed[576],seed[128],seed[2236],seed[2141],seed[696],seed[567],seed[3786],seed[1391],seed[917],seed[435],seed[313],seed[724],seed[1094],seed[1545],seed[1945],seed[1966],seed[1240],seed[1843],seed[1933],seed[3235],seed[3330],seed[1975],seed[3544],seed[2393],seed[335],seed[1453],seed[1728],seed[3301],seed[3313],seed[1173],seed[2656],seed[3957],seed[2430],seed[1570],seed[2022],seed[3024],seed[1117],seed[2247],seed[2759],seed[1497],seed[3879],seed[1855],seed[115],seed[430],seed[1078],seed[3206],seed[966],seed[3080],seed[894],seed[1585],seed[690],seed[1519],seed[518],seed[1575],seed[1556],seed[1346],seed[1214],seed[4061],seed[600],seed[4083],seed[2772],seed[2722],seed[3155],seed[424],seed[3407],seed[2638],seed[318],seed[938],seed[231],seed[781],seed[1139],seed[4009],seed[3700],seed[2540],seed[961],seed[1509],seed[3574],seed[382],seed[3520],seed[173],seed[297],seed[2483],seed[2230],seed[1192],seed[3874],seed[1398],seed[719],seed[3538],seed[1091],seed[1907],seed[1100],seed[2787],seed[3875],seed[2088],seed[2079],seed[858],seed[3469],seed[2115],seed[253],seed[536],seed[1861],seed[1761],seed[1442],seed[3279],seed[2908],seed[881],seed[3948],seed[3935],seed[2608],seed[3213],seed[3795],seed[3741],seed[3674],seed[2550],seed[3427],seed[1647],seed[2923],seed[4094],seed[429],seed[1670],seed[1491],seed[1896],seed[1439],seed[993],seed[1368],seed[2241],seed[1388],seed[2497],seed[445],seed[1464],seed[3465],seed[2127],seed[1693],seed[1521],seed[853],seed[3184],seed[2080],seed[2906],seed[11],seed[3378],seed[1134],seed[2048],seed[2380],seed[134],seed[3385],seed[2984],seed[1025],seed[1220],seed[4018],seed[3066],seed[2537],seed[1502],seed[1195]}; 
//        seed11 <= {seed[3087],seed[1951],seed[3590],seed[2376],seed[2635],seed[2218],seed[1822],seed[1923],seed[2732],seed[2860],seed[4086],seed[1029],seed[797],seed[1074],seed[2774],seed[2625],seed[338],seed[240],seed[616],seed[1283],seed[2368],seed[3039],seed[2562],seed[2865],seed[3375],seed[3057],seed[1999],seed[2116],seed[2823],seed[907],seed[856],seed[3847],seed[1514],seed[535],seed[1625],seed[2983],seed[807],seed[2746],seed[2113],seed[2094],seed[2434],seed[25],seed[1781],seed[2951],seed[1607],seed[1349],seed[1420],seed[3242],seed[3770],seed[2520],seed[1593],seed[1931],seed[1520],seed[1597],seed[3310],seed[1161],seed[813],seed[1571],seed[1254],seed[172],seed[3474],seed[2550],seed[609],seed[677],seed[2314],seed[2490],seed[3977],seed[1736],seed[3223],seed[2748],seed[1783],seed[1044],seed[2229],seed[3060],seed[3093],seed[2590],seed[3976],seed[1078],seed[1009],seed[2345],seed[1744],seed[1899],seed[2986],seed[2799],seed[660],seed[2680],seed[1488],seed[3448],seed[1250],seed[2270],seed[2644],seed[2928],seed[2016],seed[1582],seed[2864],seed[744],seed[2688],seed[66],seed[435],seed[2427],seed[2243],seed[2197],seed[1090],seed[720],seed[546],seed[689],seed[1057],seed[2668],seed[3490],seed[143],seed[2265],seed[2672],seed[2831],seed[2227],seed[2977],seed[1836],seed[1286],seed[270],seed[2666],seed[3081],seed[93],seed[1769],seed[3903],seed[787],seed[668],seed[1140],seed[750],seed[2948],seed[1155],seed[3211],seed[1208],seed[1831],seed[1542],seed[3673],seed[2740],seed[1144],seed[1911],seed[1847],seed[2246],seed[3067],seed[2226],seed[937],seed[190],seed[2964],seed[1894],seed[2463],seed[3182],seed[2884],seed[3792],seed[1401],seed[3311],seed[2881],seed[3410],seed[2543],seed[1060],seed[1065],seed[1468],seed[2082],seed[3188],seed[2849],seed[2322],seed[2030],seed[2443],seed[1082],seed[2420],seed[656],seed[265],seed[669],seed[685],seed[3080],seed[3281],seed[1369],seed[3734],seed[1383],seed[3010],seed[786],seed[3822],seed[636],seed[706],seed[3716],seed[132],seed[289],seed[2652],seed[1404],seed[2608],seed[1709],seed[3818],seed[1915],seed[432],seed[1100],seed[1224],seed[3777],seed[1813],seed[1338],seed[3220],seed[3917],seed[323],seed[2177],seed[2988],seed[2425],seed[247],seed[3268],seed[3398],seed[2313],seed[3863],seed[271],seed[124],seed[931],seed[1367],seed[2927],seed[3336],seed[407],seed[3459],seed[1977],seed[1213],seed[3186],seed[1305],seed[1067],seed[3204],seed[2115],seed[593],seed[3196],seed[2004],seed[1463],seed[2843],seed[3497],seed[3425],seed[1527],seed[905],seed[1710],seed[173],seed[2727],seed[1106],seed[2891],seed[2650],seed[2255],seed[3820],seed[3450],seed[3812],seed[625],seed[885],seed[1869],seed[2319],seed[2236],seed[886],seed[2228],seed[3793],seed[419],seed[1059],seed[178],seed[2930],seed[1551],seed[1395],seed[1350],seed[754],seed[2579],seed[1154],seed[3114],seed[2708],seed[1688],seed[153],seed[439],seed[3833],seed[3896],seed[2918],seed[1947],seed[1695],seed[332],seed[3250],seed[315],seed[1393],seed[3680],seed[1623],seed[2366],seed[1902],seed[2971],seed[2118],seed[2885],seed[3807],seed[2158],seed[48],seed[1874],seed[680],seed[227],seed[694],seed[84],seed[3049],seed[2714],seed[3688],seed[2687],seed[881],seed[3419],seed[3249],seed[3408],seed[200],seed[4014],seed[2200],seed[2621],seed[958],seed[16],seed[1330],seed[1039],seed[1760],seed[2237],seed[3644],seed[1403],seed[3523],seed[2061],seed[1515],seed[3699],seed[3533],seed[3502],seed[945],seed[2767],seed[3938],seed[2258],seed[1197],seed[2710],seed[3888],seed[1052],seed[857],seed[1231],seed[957],seed[3981],seed[2433],seed[1870],seed[1741],seed[2093],seed[2282],seed[1457],seed[3422],seed[619],seed[101],seed[0],seed[1794],seed[3233],seed[1578],seed[507],seed[1660],seed[3526],seed[1761],seed[882],seed[3573],seed[443],seed[3035],seed[2069],seed[236],seed[1469],seed[329],seed[168],seed[421],seed[1739],seed[1963],seed[1969],seed[1236],seed[3693],seed[1091],seed[3064],seed[301],seed[2701],seed[3548],seed[2691],seed[798],seed[2402],seed[2707],seed[3234],seed[2508],seed[3996],seed[513],seed[2762],seed[2492],seed[3254],seed[3559],seed[738],seed[3287],seed[2190],seed[243],seed[1827],seed[2365],seed[1173],seed[1156],seed[2855],seed[3151],seed[2092],seed[1503],seed[588],seed[1748],seed[2169],seed[2527],seed[2330],seed[461],seed[1323],seed[503],seed[1712],seed[3909],seed[1244],seed[1331],seed[2664],seed[2578],seed[836],seed[1717],seed[1664],seed[3300],seed[3374],seed[2699],seed[1662],seed[912],seed[2803],seed[3098],seed[3338],seed[795],seed[2337],seed[2937],seed[3185],seed[2396],seed[721],seed[534],seed[948],seed[708],seed[3252],seed[3208],seed[2347],seed[2769],seed[2292],seed[2859],seed[1716],seed[76],seed[966],seed[2238],seed[2995],seed[875],seed[2819],seed[2346],seed[1816],seed[1587],seed[2468],seed[2239],seed[701],seed[2060],seed[1924],seed[2012],seed[2528],seed[3030],seed[2360],seed[1158],seed[1215],seed[1528],seed[3457],seed[2309],seed[207],seed[3293],seed[3381],seed[2730],seed[3210],seed[972],seed[141],seed[3574],seed[434],seed[3106],seed[541],seed[1055],seed[3779],seed[3462],seed[3823],seed[922],seed[1363],seed[2567],seed[1177],seed[2340],seed[437],seed[41],seed[1989],seed[902],seed[691],seed[2025],seed[3386],seed[2268],seed[455],seed[2382],seed[2580],seed[2168],seed[1202],seed[206],seed[898],seed[108],seed[852],seed[1324],seed[3889],seed[1719],seed[194],seed[2195],seed[3238],seed[2599],seed[3536],seed[122],seed[1497],seed[3356],seed[2614],seed[2934],seed[3253],seed[2047],seed[2291],seed[220],seed[2601],seed[4030],seed[1512],seed[4059],seed[2645],seed[5],seed[1807],seed[2775],seed[3984],seed[3277],seed[2872],seed[3218],seed[468],seed[1507],seed[3148],seed[341],seed[2355],seed[1178],seed[2682],seed[1088],seed[878],seed[3668],seed[1408],seed[2096],seed[2690],seed[2628],seed[3513],seed[1934],seed[3146],seed[2811],seed[2956],seed[1269],seed[1170],seed[1801],seed[1113],seed[2377],seed[1960],seed[3529],seed[3470],seed[1336],seed[1282],seed[3487],seed[556],seed[3028],seed[831],seed[695],seed[1653],seed[648],seed[217],seed[3610],seed[2828],seed[43],seed[339],seed[768],seed[3364],seed[1583],seed[2479],seed[2585],seed[3525],seed[3906],seed[318],seed[1255],seed[3550],seed[3138],seed[26],seed[2077],seed[2009],seed[1412],seed[3388],seed[2893],seed[3316],seed[2801],seed[2406],seed[2835],seed[523],seed[2968],seed[3508],seed[2279],seed[2572],seed[1204],seed[2136],seed[1610],seed[1038],seed[3290],seed[994],seed[1217],seed[3510],seed[3436],seed[1428],seed[911],seed[3011],seed[2633],seed[3911],seed[3446],seed[2328],seed[1212],seed[1049],seed[1141],seed[1838],seed[3702],seed[3578],seed[3475],seed[2686],seed[4068],seed[1810],seed[110],seed[1536],seed[3382],seed[568],seed[2189],seed[1697],seed[2401],seed[2233],seed[2250],seed[672],seed[1480],seed[3163],seed[1313],seed[1658],seed[1157],seed[3541],seed[801],seed[575],seed[4026],seed[2700],seed[773],seed[557],seed[973],seed[377],seed[1132],seed[397],seed[819],seed[4043],seed[1203],seed[2208],seed[2657],seed[1600],seed[3484],seed[1419],seed[152],seed[245],seed[3278],seed[2674],seed[2491],seed[2219],seed[2153],seed[55],seed[1601],seed[3391],seed[3222],seed[3625],seed[2648],seed[2742],seed[3308],seed[2834],seed[412],seed[3275],seed[3582],seed[3442],seed[1855],seed[3692],seed[3885],seed[1133],seed[743],seed[1853],seed[942],seed[3133],seed[3841],seed[2901],seed[1438],seed[3379],seed[3845],seed[2825],seed[29],seed[848],seed[3443],seed[2619],seed[2387],seed[1421],seed[1517],seed[510],seed[3890],seed[325],seed[985],seed[2119],seed[3628],seed[1817],seed[1056],seed[1168],seed[2217],seed[3344],seed[330],seed[46],seed[757],seed[401],seed[1939],seed[2157],seed[361],seed[1406],seed[1701],seed[1698],seed[2424],seed[4007],seed[698],seed[3198],seed[4058],seed[3961],seed[1198],seed[2352],seed[3922],seed[3272],seed[3972],seed[1543],seed[1700],seed[3165],seed[3875],seed[2139],seed[969],seed[3740],seed[2059],seed[2594],seed[1477],seed[3848],seed[1071],seed[1627],seed[4063],seed[2498],seed[1879],seed[3763],seed[1998],seed[2669],seed[1342],seed[1117],seed[2416],seed[250],seed[2461],seed[293],seed[3018],seed[3866],seed[1092],seed[2404],seed[3825],seed[1859],seed[224],seed[612],seed[747],seed[4018],seed[335],seed[1549],seed[1928],seed[1353],seed[3140],seed[3147],seed[884],seed[2904],seed[3775],seed[4047],seed[149],seed[452],seed[2781],seed[1301],seed[2362],seed[1704],seed[3506],seed[3321],seed[1464],seed[955],seed[967],seed[3879],seed[2902],seed[3636],seed[2123],seed[1222],seed[4019],seed[1162],seed[3561],seed[2386],seed[1667],seed[1793],seed[3608],seed[1680],seed[3413],seed[2180],seed[1247],seed[133],seed[587],seed[1945],seed[13],seed[2676],seed[2571],seed[2028],seed[815],seed[2378],seed[2138],seed[1315],seed[3320],seed[1965],seed[765],seed[2761],seed[3751],seed[904],seed[1436],seed[1973],seed[1297],seed[779],seed[1192],seed[258],seed[482],seed[2288],seed[628],seed[2205],seed[2895],seed[1278],seed[1196],seed[3135],seed[1509],seed[286],seed[563],seed[3919],seed[1252],seed[1656],seed[1304],seed[1339],seed[59],seed[3167],seed[756],seed[1502],seed[572],seed[722],seed[2379],seed[1239],seed[3373],seed[2867],seed[2494],seed[1575],seed[1399],seed[2369],seed[2220],seed[724],seed[1312],seed[1351],seed[3784],seed[2080],seed[538],seed[3161],seed[1833],seed[3748],seed[1111],seed[209],seed[2310],seed[2040],seed[3685],seed[3362],seed[488],seed[2500],seed[2182],seed[1755],seed[959],seed[2400],seed[1063],seed[415],seed[2752],seed[1628],seed[204],seed[3988],seed[591],seed[3819],seed[2763],seed[2114],seed[2445],seed[2336],seed[1216],seed[3332],seed[2624],seed[1424],seed[203],seed[371],seed[1279],seed[3665],seed[639],seed[3267],seed[1040],seed[277],seed[3957],seed[617],seed[1830],seed[2364],seed[1839],seed[4006],seed[2496],seed[1579],seed[3766],seed[2058],seed[979],seed[1182],seed[1249],seed[2531],seed[1335],seed[3318],seed[2980],seed[4055],seed[584],seed[1572],seed[3724],seed[2050],seed[2423],seed[1577],seed[3342],seed[3966],seed[4090],seed[3058],seed[2470],seed[2792],seed[734],seed[991],seed[2514],seed[586],seed[296],seed[2609],seed[3444],seed[2501],seed[1584],seed[1455],seed[2861],seed[3472],seed[2512],seed[350],seed[2539],seed[2641],seed[1373],seed[1861],seed[3681],seed[1083],seed[3645],seed[242],seed[3224],seed[3517],seed[2517],seed[1409],seed[281],seed[1491],seed[3024],seed[462],seed[2341],seed[1532],seed[2737],seed[1261],seed[3677],seed[626],seed[2043],seed[279],seed[1670],seed[3746],seed[1445],seed[543],seed[3191],seed[316],seed[1745],seed[598],seed[3756],seed[1073],seed[2909],seed[1903],seed[1325],seed[3121],seed[2804],seed[2758],seed[897],seed[302],seed[1955],seed[1362],seed[599],seed[3285],seed[15],seed[3447],seed[3619],seed[2155],seed[2034],seed[3044],seed[1019],seed[19],seed[3799],seed[771],seed[72],seed[1030],seed[1461],seed[566],seed[3393],seed[2171],seed[3893],seed[2906],seed[2681],seed[1268],seed[4085],seed[3181],seed[2485],seed[38],seed[2176],seed[1416],seed[3117],seed[711],seed[3205],seed[3542],seed[3059],seed[2592],seed[1322],seed[2962],seed[365],seed[1865],seed[1636],seed[1620],seed[2894],seed[3498],seed[1103],seed[60],seed[2754],seed[3209],seed[1237],seed[478],seed[2502],seed[3183],seed[1129],seed[3515],seed[363],seed[3620],seed[870],seed[3461],seed[1518],seed[1771],seed[638],seed[3778],seed[3020],seed[1715],seed[834],seed[2163],seed[3760],seed[3296],seed[675],seed[3733],seed[950],seed[2534],seed[2837],seed[2407],seed[2221],seed[8],seed[3331],seed[3309],seed[3108],seed[2278],seed[1242],seed[627],seed[3495],seed[1529],seed[849],seed[3325],seed[3654],seed[3271],seed[4020],seed[2982],seed[1631],seed[1863],seed[2194],seed[1886],seed[3789],seed[1702],seed[233],seed[3232],seed[1824],seed[2390],seed[1589],seed[883],seed[1504],seed[1022],seed[491],seed[234],seed[2908],seed[2515],seed[3759],seed[2342],seed[2991],seed[2356],seed[2032],seed[2544],seed[1691],seed[1214],seed[3951],seed[2844],seed[3174],seed[2324],seed[1265],seed[3967],seed[2411],seed[1940],seed[1634],seed[117],seed[1565],seed[1025],seed[1172],seed[1720],seed[2274],seed[3660],seed[2299],seed[895],seed[2802],seed[3125],seed[3821],seed[1333],seed[1825],seed[624],seed[3006],seed[3797],seed[1291],seed[2551],seed[492],seed[411],seed[1318],seed[2576],seed[3736],seed[2394],seed[3496],seed[929],seed[903],seed[274],seed[3745],seed[2399],seed[3642],seed[358],seed[2188],seed[1981],seed[3894],seed[120],seed[1788],seed[257],seed[2117],seed[2665],seed[67],seed[3708],seed[1867],seed[3110],seed[3786],seed[2606],seed[601],seed[3123],seed[1506],seed[3492],seed[1273],seed[3883],seed[2888],seed[3068],seed[1950],seed[2482],seed[3377],seed[3101],seed[2890],seed[3257],seed[3678],seed[936],seed[3588],seed[2143],seed[4001],seed[1987],seed[2677],seed[450],seed[2555],seed[2022],seed[3920],seed[683],seed[1659],seed[2466],seed[2945],seed[533],seed[1522],seed[654],seed[2134],seed[3430],seed[2879],seed[2979],seed[3458],seed[1516],seed[865],seed[174],seed[1189],seed[3322],seed[673],seed[1699],seed[632],seed[550],seed[3276],seed[3768],seed[106],seed[820],seed[2430],seed[1780],seed[2041],seed[116],seed[3900],seed[410],seed[2137],seed[2753],seed[2751],seed[9],seed[163],seed[1472],seed[2006],seed[2653],seed[3960],seed[304],seed[288],seed[841],seed[3750],seed[611],seed[551],seed[3511],seed[1602],seed[2846],seed[4060],seed[3399],seed[33],seed[2790],seed[1240],seed[2505],seed[3916],seed[3004],seed[2241],seed[3732],seed[324],seed[1980],seed[811],seed[2773],seed[1875],seed[613],seed[582],seed[3134],seed[1718],seed[3184],seed[1734],seed[3571],seed[1102],seed[3107],seed[536],seed[2726],seed[2974],seed[2807],seed[1731],seed[581],seed[2993],seed[2211],seed[714],seed[3586],seed[2214],seed[334],seed[1035],seed[728],seed[2325],seed[2405],seed[2911],seed[3500],seed[1724],seed[1918],seed[571],seed[1145],seed[3111],seed[1459],seed[3397],seed[405],seed[2320],seed[3555],seed[901],seed[3126],seed[956],seed[1791],seed[2910],seed[2283],seed[2141],seed[3481],seed[3292],seed[3017],seed[4037],seed[1893],seed[2970],seed[112],seed[1892],seed[1941],seed[2581],seed[3159],seed[1443],seed[4061],seed[80],seed[2583],seed[1654],seed[3664],seed[1535],seed[322],seed[3061],seed[3479],seed[604],seed[3537],seed[438],seed[2734],seed[1176],seed[4067],seed[3927],seed[3880],seed[1066],seed[3274],seed[1513],seed[3964],seed[1064],seed[2230],seed[1042],seed[2719],seed[2586],seed[1200],seed[3622],seed[2079],seed[2656],seed[1851],seed[1606],seed[791],seed[4070],seed[840],seed[4003],seed[3728],seed[2179],seed[1316],seed[1835],seed[2874],seed[2617],seed[2454],seed[2263],seed[352],seed[1233],seed[2375],seed[2838],seed[2965],seed[1046],seed[3266],seed[1953],seed[818],seed[2822],seed[63],seed[540],seed[858],seed[346],seed[781],seed[208],seed[1364],seed[425],seed[3790],seed[2703],seed[3130],seed[388],seed[3593],seed[780],seed[3306],seed[3008],seed[2866],seed[1006],seed[2472],seed[2088],seed[923],seed[2172],seed[3164],seed[3902],seed[184],seed[2304],seed[487],seed[3783],seed[483],seed[971],seed[2484],seed[3547],seed[1540],seed[1377],seed[1806],seed[305],seed[31],seed[2836],seed[2308],seed[3684],seed[1763],seed[3007],seed[269],seed[2152],seed[1084],seed[3414],seed[2778],seed[3721],seed[1622],seed[2671],seed[2743],seed[1328],seed[1531],seed[195],seed[3023],seed[453],seed[248],seed[3549],seed[2344],seed[2526],seed[2202],seed[3371],seed[2768],seed[2286],seed[1034],seed[1195],seed[2728],seed[1795],seed[3473],seed[2223],seed[3899],seed[2622],seed[3323],seed[1206],seed[3137],seed[2694],seed[140],seed[938],seed[4044],seed[2765],seed[740],seed[3389],seed[3225],seed[1276],seed[2588],seed[376],seed[480],seed[1792],seed[87],seed[2244],seed[1302],seed[845],seed[1184],seed[463],seed[3962],seed[1394],seed[1842],seed[4084],seed[62],seed[1677],seed[3904],seed[254],seed[386],seed[4074],seed[3709],seed[327],seed[3915],seed[57],seed[761],seed[3602],seed[2389],seed[1614],seed[40],seed[3861],seed[1845],seed[3801],seed[3539],seed[3910],seed[846],seed[860],seed[3752],seed[157],seed[71],seed[264],seed[3887],seed[879],seed[2791],seed[369],seed[3580],seed[3767],seed[1686],seed[23],seed[1451],seed[3772],seed[1434],seed[2412],seed[3143],seed[3019],seed[1804],seed[2135],seed[299],seed[2480],seed[3924],seed[981],seed[690],seed[1905],seed[1674],seed[2207],seed[3975],seed[1714],seed[953],seed[2145],seed[3201],seed[3862],seed[3959],seed[640],seed[298],seed[3109],seed[256],seed[3715],seed[1519],seed[2827],seed[1889],seed[3992],seed[3],seed[24],seed[866],seed[3226],seed[1984],seed[1016],seed[987],seed[3969],seed[3579],seed[3269],seed[1450],seed[105],seed[1109],seed[3616],seed[3097],seed[1815],seed[130],seed[2736],seed[4029],seed[800],seed[441],seed[916],seed[2005],seed[1913],seed[2613],seed[589],seed[1346],seed[996],seed[3273],seed[3365],seed[1124],seed[2563],seed[1169],seed[592],seed[3613],seed[578],seed[1258],seed[1872],seed[1558],seed[2095],seed[2558],seed[3738],seed[394],seed[862],seed[2109],seed[1388],seed[4032],seed[1385],seed[1199],seed[3735],seed[1372],seed[2772],seed[1900],seed[1541],seed[3380],seed[2738],seed[1723],seed[2306],seed[662],seed[1562],seed[2224],seed[3353],seed[2955],seed[3084],seed[1048],seed[2293],seed[716],seed[2718],seed[2545],seed[700],seed[2771],seed[603],seed[3634],seed[995],seed[1611],seed[3546],seed[2146],seed[2165],seed[1221],seed[2075],seed[2932],seed[3319],seed[2410],seed[3394],seed[420],seed[3742],seed[175],seed[3343],seed[736],seed[2462],seed[1164],seed[4049],seed[3597],seed[2056],seed[3015],seed[192],seed[1422],seed[3095],seed[2642],seed[2994],seed[3757],seed[37],seed[2240],seed[3871],seed[1390],seed[2072],seed[4089],seed[4028],seed[3070],seed[1024],seed[4094],seed[1511],seed[3519],seed[2729],seed[1460],seed[2961],seed[3054],seed[1895],seed[2770],seed[3217],seed[287],seed[2784],seed[1678],seed[3596],seed[876],seed[2915],seed[2002],seed[131],seed[1959],seed[460],seed[3557],seed[2739],seed[2854],seed[2083],seed[2478],seed[2654],seed[310],seed[1896],seed[3970],seed[692],seed[1290],seed[827],seed[2914],seed[3648],seed[3706],seed[3698],seed[3753],seed[1742],seed[2196],seed[121],seed[835],seed[775],seed[2535],seed[3466],seed[2851],seed[686],seed[3844],seed[177],seed[2840],seed[4065],seed[1020],seed[3810],seed[1707],seed[1128],seed[2936],seed[2024],seed[1938],seed[3357],seed[1689],seed[2298],seed[1966],seed[2800],seed[717],seed[3946],seed[3552],seed[2052],seed[1823],seed[1452],seed[424],seed[645],seed[1355],seed[788],seed[50],seed[171],seed[3100],seed[2327],seed[2570],seed[445],seed[490],seed[3166],seed[799],seed[1160],seed[147],seed[682],seed[1287],seed[1292],seed[447],seed[1310],seed[366],seed[782],seed[1849],seed[2252],seed[4015],seed[2873],seed[3505],seed[3929],seed[2667],seed[3605],seed[210],seed[56],seed[888],seed[252],seed[529],seed[674],seed[3538],seed[1776],seed[212],seed[1566],seed[3626],seed[2921],seed[2805],seed[241],seed[73],seed[356],seed[349],seed[2939],seed[2826],seed[553],seed[3348],seed[1777],seed[3301],seed[2105],seed[1501],seed[3088],seed[3305],seed[3485],seed[2992],seed[3575],seed[2184],seed[2388],seed[2573],seed[393],seed[1238],seed[3788],seed[3884],seed[3993],seed[3177],seed[3075],seed[3445],seed[3858],seed[1877],seed[594],seed[3621],seed[2003],seed[2107],seed[2036],seed[3467],seed[3132],seed[505],seed[4093],seed[837],seed[558],seed[2102],seed[3477],seed[3944],seed[1770],seed[499],seed[3045],seed[2483],seed[1733],seed[1829],seed[1475],seed[3898],seed[2091],seed[1314],seed[36],seed[2133],seed[3424],seed[2733],seed[68],seed[528],seed[947],seed[3040],seed[3429],seed[1661],seed[2756],seed[3982],seed[30],seed[1473],seed[1616],seed[774],seed[1946],seed[3435],seed[1079],seed[1919],seed[2090],seed[2919],seed[278],seed[1007],seed[684],seed[1901],seed[3565],seed[3014],seed[1643],seed[3791],seed[1843],seed[2029],seed[2725],seed[474],seed[968],seed[99],seed[2000],seed[90],seed[1326],seed[735],seed[2267],seed[1442],seed[2206],seed[2941],seed[2582],seed[1123],seed[2186],seed[778],seed[642],seed[385],seed[2847],seed[1922],seed[235],seed[2457],seed[1440],seed[2301],seed[225],seed[3284],seed[2552],seed[1560],seed[3874],seed[403],seed[17],seed[2048],seed[1487],seed[2812],seed[926],seed[1706],seed[1858],seed[928],seed[2824],seed[198],seed[2780],seed[1075],seed[231],seed[211],seed[3953],seed[3086],seed[2522],seed[3599],seed[951],seed[542],seed[268],seed[3417],seed[833],seed[2931],seed[3703],seed[158],seed[381],seed[4048],seed[21],seed[473],seed[2486],seed[3094],seed[3501],seed[3175],seed[2063],seed[1226],seed[637],seed[1649],seed[4054],seed[2487],seed[2357],seed[2277],seed[1604],seed[2385],seed[3947],seed[1142],seed[2380],seed[100],seed[2110],seed[3631],seed[699],seed[4009],seed[1288],seed[1370],seed[1917],seed[1613],seed[308],seed[3646],seed[185],seed[1332],seed[1635],seed[1219],seed[1975],seed[1995],seed[230],seed[1942],seed[939],seed[3170],seed[3998],seed[671],seed[3794],seed[1873],seed[2549],seed[1568],seed[3345],seed[4010],seed[2816],seed[1642],seed[3295],seed[3923],seed[3199],seed[2130],seed[493],seed[484],seed[3187],seed[2162],seed[564],seed[1876],seed[2720],seed[1651],seed[3326],seed[3216],seed[2721],seed[2348],seed[199],seed[237],seed[11],seed[1340],seed[418],seed[2913],seed[4004],seed[696],seed[896],seed[426],seed[3744],seed[454],seed[917],seed[1054],seed[2010],seed[1799],seed[3531],seed[1929],seed[54],seed[2448],seed[1131],seed[605],seed[580],seed[1805],seed[3643],seed[577],seed[1274],seed[1345],seed[3989],seed[2593],seed[3630],seed[3564],seed[3554],seed[3999],seed[176],seed[78],seed[3667],seed[1703],seed[3925],seed[2132],seed[1347],seed[954],seed[2821],seed[4005],seed[3179],seed[2326],seed[3178],seed[34],seed[1967],seed[3297],seed[164],seed[746],seed[359],seed[3815],seed[2493],seed[1094],seed[1976],seed[3609],seed[1721],seed[357],seed[4038],seed[3160],seed[3193],seed[3892],seed[2111],seed[2958],seed[2875],seed[3259],seed[1391],seed[812],seed[2541],seed[2422],seed[2598],seed[2519],seed[687],seed[3263],seed[576],seed[1914],seed[440],seed[1118],seed[282],seed[317],seed[1790],seed[2343],seed[2722],seed[3651],seed[3085],seed[408],seed[1045],seed[3158],seed[1309],seed[3504],seed[2981],seed[3935],seed[221],seed[732],seed[518],seed[935],seed[3033],seed[3905],seed[3482],seed[2297],seed[1537],seed[2311],seed[1003],seed[1293],seed[3842],seed[1115],seed[3516],seed[2011],seed[1961],seed[597],seed[3229],seed[2391],seed[545],seed[2154],seed[2068],seed[3346],seed[2247],seed[1474],seed[2692],seed[1585],seed[2333],seed[2705],seed[1814],seed[3456],seed[1259],seed[2757],seed[650],seed[88],seed[2216],seed[396],seed[1526],seed[3197],seed[952],seed[4017],seed[1467],seed[2307],seed[2697],seed[20],seed[3816],seed[2521],seed[2354],seed[2349],seed[2264],seed[3053],seed[2950],seed[1486],seed[3120],seed[2167],seed[1068],seed[4045],seed[517],seed[2525],seed[1187],seed[1605],seed[2149],seed[2985],seed[806],seed[1281],seed[2103],seed[2611],seed[3583],seed[2323],seed[3401],seed[364],seed[579],seed[1190],seed[2712],seed[1997],seed[755],seed[1750],seed[69],seed[370],seed[697],seed[3945],seed[3682],seed[569],seed[1878],seed[3455],seed[1081],seed[3983],seed[1228],seed[2225],seed[2023],seed[688],seed[4064],seed[565],seed[3776],seed[253],seed[4025],seed[2131],seed[1303],seed[1725],seed[1523],seed[3612],seed[520],seed[2600],seed[817],seed[3129],seed[2312],seed[678],seed[863],seed[1949],seed[1818],seed[659],seed[368],seed[3432],seed[512],seed[1621],seed[3584],seed[2536],seed[1789],seed[2395],seed[3215],seed[404],seed[3029],seed[2201],seed[1772],seed[306],seed[2474],seed[2151],seed[3627],seed[1671],seed[1225],seed[3113],seed[670],seed[3876],seed[391],seed[667],seed[2446],seed[1398],seed[4091],seed[2066],seed[760],seed[552],seed[2627],seed[2044],seed[2419],seed[3921],seed[1307],seed[3878],seed[2317],seed[267],seed[918],seed[1134],seed[1116],seed[1569],seed[2035],seed[326],seed[1396],seed[3831],seed[1483],seed[3869],seed[3840],seed[1666],seed[871],seed[2749],seed[1193],seed[1402],seed[3384],seed[2129],seed[2537],seed[126],seed[223],seed[2042],seed[3050],seed[10],seed[877],seed[851],seed[295],seed[2510],seed[2475],seed[867],seed[2833],seed[2261],seed[154],seed[4053],seed[949],seed[1751],seed[766],seed[3036],seed[3641],seed[1880],seed[1361],seed[3737],seed[3963],seed[3065],seed[2695],seed[531],seed[2513],seed[1758],seed[2335],seed[2099],seed[1599],seed[2516],seed[2876],seed[3572],seed[2880],seed[1061],seed[1834],seed[749],seed[653],seed[2820],seed[1137],seed[2440],seed[502],seed[3679],seed[1740],seed[2212],seed[1496],seed[1076],seed[839],seed[2946],seed[3051],seed[3800],seed[934],seed[2848],seed[664],seed[1548],seed[1920],seed[514],seed[2696],seed[3202],seed[2465],seed[1538],seed[1080],seed[2124],seed[390],seed[1673],seed[1356],seed[1550],seed[4039],seed[1580],seed[494],seed[2886],seed[1738],seed[1485],seed[1809],seed[789],seed[2358],seed[2810],seed[854],seed[465],seed[1767],seed[2912],seed[2796],seed[2612],seed[1209],seed[1433],seed[1058],seed[1146],seed[2561],seed[2639],seed[1023],seed[629],seed[150],seed[2101],seed[3241],seed[1907],seed[2683],seed[3071],seed[3207],seed[2019],seed[2923],seed[3280],seed[3037],seed[983],seed[1185],seed[3089],seed[899],seed[3524],seed[1037],seed[161],seed[1525],seed[3918],seed[2017],seed[993],seed[2222],seed[111],seed[179],seed[2020],seed[3031],seed[615],seed[1754],seed[2026],seed[1267],seed[2271],seed[219],seed[2907],seed[3696],seed[3867],seed[3663],seed[2530],seed[98],seed[2269],seed[2495],seed[2862],seed[707],seed[2659],seed[3615],seed[181],seed[442],seed[1898],seed[1150],seed[1624],seed[64],seed[1684],seed[2591],seed[1775],seed[3676],seed[3873],seed[1337],seed[340],seed[3282],seed[3073],seed[2776],seed[537],seed[413],seed[2213],seed[1985],seed[3079],seed[2021],seed[2147],seed[1581],seed[1676],seed[906],seed[337],seed[880],seed[94],seed[3337],seed[1234],seed[3958],seed[2903],seed[1968],seed[3623],seed[162],seed[1832],seed[3830],seed[2262],seed[3192],seed[1639],seed[1354],seed[1375],seed[3769],seed[3639],seed[777],seed[3270],seed[2808],seed[2159],seed[1533],seed[1223],seed[259],seed[2996],seed[3152],seed[2782],seed[1557],seed[2741],seed[3145],seed[65],seed[3859],seed[351],seed[3043],seed[205],seed[1021],seed[1295],seed[1904],seed[2787],seed[3055],seed[1435],seed[3581],seed[2603],seed[3324],seed[2938],seed[988],seed[4042],seed[3335],seed[3881],seed[3624],seed[3758],seed[1490],seed[2086],seed[1005],seed[1425],seed[1728],seed[3534],seed[1389],seed[61],seed[2361],seed[3591],seed[3453],seed[2100],seed[2421],seed[3312],seed[372],seed[727],seed[1826],seed[2646],seed[2473],seed[3489],seed[2174],seed[47],seed[1341],seed[1713],seed[4051],seed[665],seed[2070],seed[486],seed[1881],seed[792],seed[965],seed[2713],seed[3955],seed[1050],seed[2497],seed[436],seed[2334],seed[1018],seed[2393],seed[2458],seed[255],seed[3601],seed[3979],seed[2518],seed[753],seed[284],seed[4035],seed[3544],seed[448],seed[821],seed[3025],seed[509],seed[1366],seed[1494],seed[417],seed[3483],seed[3817],seed[427],seed[618],seed[3299],seed[1800],seed[374],seed[1028],seed[320],seed[1479],seed[631],seed[655],seed[1382],seed[3700],seed[280],seed[853],seed[28],seed[1499],seed[1640],seed[893],seed[1685],seed[3978],seed[1521],seed[1194],seed[1837],seed[1426],seed[784],seed[1218],seed[1343],seed[2128],seed[2367],seed[3153],seed[3291],seed[3072],seed[3705],seed[2899],seed[1737],seed[3460],seed[229],seed[2717],seed[3009],seed[2455],seed[2856],seed[1013],seed[2850],seed[2084],seed[2640],seed[2998],seed[2973],seed[977],seed[2256],seed[495],seed[1498],seed[1149],seed[960],seed[770],seed[1031],seed[3361],seed[389],seed[3122],seed[1983],seed[251],seed[3826],seed[2284],seed[2183],seed[1693],seed[4],seed[314],seed[829],seed[1381],seed[1598],seed[3206],seed[1120],seed[3614],seed[2467],seed[1026],seed[1570],seed[414],seed[567],seed[1047],seed[3387],seed[2046],seed[1386],seed[525],seed[2702],seed[2148],seed[3814],seed[1348],seed[2632],seed[354],seed[2935],seed[676],seed[2234],seed[3131],seed[1906],seed[3604],seed[1812],seed[4072],seed[2623],seed[2809],seed[3687],seed[3251],seed[1476],seed[187],seed[3118],seed[3697],seed[718],seed[925],seed[1112],seed[1927],seed[963],seed[3368],seed[2418],seed[1668],seed[1840],seed[3811],seed[2967],seed[3156],seed[1500],seed[2477],seed[4022],seed[3235],seed[872],seed[526],seed[2359],seed[2429],seed[3367],seed[772],seed[530],seed[2924],seed[816],seed[574],seed[3839],seed[1746],seed[1344],seed[1596],seed[3303],seed[661],seed[3330],seed[2877],seed[1441],seed[793],seed[3013],seed[830],seed[2015],seed[2232],seed[290],seed[3162],seed[710],seed[3418],seed[2013],seed[726],seed[294],seed[2673],seed[3710],seed[2715],seed[3124],seed[1785],seed[3294],seed[1179],seed[719],seed[3228],seed[3527],seed[409],seed[3240],seed[1300],seed[2332],seed[997],seed[74],seed[3434],seed[2456],seed[2795],seed[3358],seed[1165],seed[2081],seed[3077],seed[261],seed[962],seed[497],seed[3265],seed[2607],seed[910],seed[1053],seed[2417],seed[123],seed[2698],seed[2315],seed[1629],seed[3403],seed[213],seed[226],seed[713],seed[1368],seed[560],seed[1387],seed[1456],seed[3658],seed[2731],seed[3701],seed[2442],seed[382],seed[1730],seed[2589],seed[3244],seed[992],seed[1682],seed[3933],seed[850],seed[1360],seed[2871],seed[3834],seed[3870],seed[3649],seed[3857],seed[1321],seed[2481],seed[3617],seed[3376],seed[1756],seed[138],seed[3493],seed[2660],seed[2560],seed[3592],seed[2538],seed[1122],seed[3854],seed[4000],seed[1308],seed[1595],seed[3528],seed[1256],seed[331],seed[3115],seed[3606],seed[2173],seed[1862],seed[4095],seed[2089],seed[3942],seed[2533],seed[2777],seed[1732],seed[3359],seed[1552],seed[3069],seed[3940],seed[1033],seed[51],seed[2464],seed[1787],seed[3354],seed[519],seed[3836],seed[606],seed[367],seed[1207],seed[2053],seed[1856],seed[3426],seed[1774],seed[1972],seed[1753],seed[3214],seed[3828],seed[693],seed[908],seed[1888],seed[3675],seed[873],seed[3339],seed[3105],seed[741],seed[489],seed[2381],seed[2595],seed[3363],seed[1],seed[4040],seed[3407],seed[3743],seed[4075],seed[3427],seed[3633],seed[3454],seed[602],seed[643],seed[3587],seed[2450],seed[1235],seed[501],seed[1495],seed[1743],seed[197],seed[2447],seed[1069],seed[3856],seed[3022],seed[2126],seed[3333],seed[1645],seed[2989],seed[4077],seed[3670],seed[946],seed[469],seed[428],seed[737],seed[1726],seed[2832],seed[1493],seed[559],seed[2351],seed[2295],seed[3149],seed[3635],seed[3686],seed[2916],seed[1272],seed[1334],seed[2897],seed[2815],seed[1964],seed[2414],seed[3431],seed[169],seed[1296],seed[1908],seed[2779],seed[3991],seed[2630],seed[2735],seed[3607],seed[3829],seed[842],seed[1930],seed[3808],seed[3535],seed[3749],seed[2038],seed[742],seed[1077],seed[2987],seed[767],seed[3005],seed[986],seed[3136],seed[113],seed[3260],seed[2529],seed[2018],seed[1107],seed[3180],seed[3027],seed[2372],seed[3707],seed[3913],seed[3914],seed[3827],seed[4062],seed[1166],seed[472],seed[1163],seed[3930],seed[2556],seed[344],seed[500],seed[430],seed[360],seed[2905],seed[2409],seed[2532],seed[874],seed[3046],seed[3503],seed[1125],seed[4041],seed[964],seed[2403],seed[620],seed[2187],seed[725],seed[2511],seed[3416],seed[583],seed[58],seed[3347],seed[1482],seed[3433],seed[1974],seed[1484],seed[3780],seed[238],seed[2542],seed[1201],seed[3860],seed[2062],seed[703],seed[1802],seed[244],seed[943],seed[1379],seed[2209],seed[2441],seed[855],seed[1808],seed[466],seed[218],seed[3279],seed[2453],seed[2087],seed[1138],seed[2296],seed[1608],seed[2127],seed[1937],seed[2120],seed[2643],seed[475],seed[3567],seed[1284],seed[1933],seed[2249],seed[1594],seed[1996],seed[193],seed[2275],seed[1220],seed[347],seed[1555],seed[3518],seed[3562],seed[608],seed[2305],seed[824],seed[2723],seed[2892],seed[1576],seed[832],seed[136],seed[375],seed[823],seed[1979],seed[186],seed[1015],seed[3203],seed[109],seed[1641],seed[941],seed[802],seed[155],seed[914],seed[1971],seed[52],seed[3091],seed[456],seed[3719],seed[2689],seed[1764],seed[532],seed[311],seed[554],seed[3994],seed[894],seed[3421],seed[3420],seed[2917],seed[3712],seed[196],seed[3928],seed[3809],seed[2870],seed[3247],seed[3986],seed[160],seed[1264],seed[3603],seed[1243],seed[887],seed[890],seed[128],seed[1263],seed[2788],seed[3973],seed[2428],seed[2944],seed[1119],seed[3486],seed[3001],seed[3314],seed[1289],seed[915],seed[2574],seed[2242],seed[1567],seed[1615],seed[2300],seed[2098],seed[859],seed[82],seed[433],seed[2488],seed[561],seed[1637],seed[3449],seed[214],seed[3837],seed[3666],seed[1374],seed[3764],seed[614],seed[2755],seed[2122],seed[479],seed[808],seed[1657],seed[3931],seed[2266],seed[2631],seed[2259],seed[3150],seed[3480],seed[3852],seed[3689],seed[2553],seed[1087],seed[328],seed[635],seed[2959],seed[1821],seed[2460],seed[745],seed[1988],seed[2814],seed[1405],seed[3230],seed[406],seed[2947],seed[647],seed[1683],seed[3127],seed[292],seed[3315],seed[395],seed[127],seed[2798],seed[1803],seed[1708],seed[12],seed[809],seed[3835],seed[1786],seed[3169],seed[1854],seed[1883],seed[2104],seed[1935],seed[1530],seed[3730],seed[1962],seed[3901],seed[4023],seed[2818],seed[142],seed[3585],seed[3514],seed[429],seed[555],seed[1104],seed[3385],seed[610],seed[1481],seed[1175],seed[3369],seed[1210],seed[2185],seed[2384],seed[4050],seed[89],seed[97],seed[3674],seed[527],seed[1152],seed[3441],seed[1257],seed[2602],seed[1086],seed[2557],seed[1864],seed[1779],seed[151],seed[3632],seed[2675],seed[3509],seed[342],seed[39],seed[658],seed[1097],seed[2064],seed[2074],seed[77],seed[3438],seed[2651],seed[336],seed[3711],seed[1958],seed[146],seed[400],seed[1089],seed[2193],seed[1446],seed[2051],seed[2008],seed[1127],seed[1151],seed[42],seed[3761],seed[4013],seed[2786],seed[3262],seed[1705],seed[4071],seed[731],seed[1099],seed[1191],seed[348],seed[2637],seed[573],seed[2957],seed[2371],seed[2963],seed[3722],seed[2204],seed[139],seed[759],seed[2662],seed[3556],seed[215],seed[2353],seed[1266],seed[1384],seed[1130],seed[4027],seed[621],seed[3714],seed[3655],seed[657],seed[1954],seed[353],seed[1638],seed[2142],seed[3392],seed[3112],seed[3016],seed[2031],seed[3428],seed[3908],seed[4031],seed[4081],seed[1432],seed[3200],seed[1148],seed[2503],seed[1271],seed[2476],seed[3803],seed[3650],seed[590],seed[3465],seed[864],seed[3038],seed[2459],seed[1153],seed[2285],seed[2439],seed[2615],seed[3595],seed[2260],seed[81],seed[1466],seed[630],seed[300],seed[3056],seed[2817],seed[2280],seed[159],seed[3494],seed[2469],seed[3782],seed[1765],seed[3237],seed[2565],seed[932],seed[805],seed[1553],seed[3003],seed[3302],seed[2408],seed[733],seed[1458],seed[3941],seed[3404],seed[3865],seed[2604],seed[764],seed[2281],seed[457],seed[3173],seed[3741],seed[95],seed[3212],seed[2852],seed[3390],seed[2597],seed[3600],seed[3838],seed[1675],seed[2922],seed[3372],seed[2125],seed[1471],seed[321],seed[1010],seed[2071],seed[652],seed[1992],seed[1603],seed[1650],seed[1327],seed[1357],seed[392],seed[1085],seed[2289],seed[1564],seed[398],seed[423],seed[431],seed[1711],seed[1311],seed[1147],seed[4033],seed[1912],seed[1563],seed[144],seed[44],seed[103],seed[2150],seed[3569],seed[3261],seed[3154],seed[3116],seed[2661],seed[521],seed[2057],seed[3488],seed[3798],seed[1952],seed[4080],seed[3440],seed[3577],seed[1245],seed[3720],seed[646],seed[3553],seed[1665],seed[1043],seed[1262],seed[1647],seed[2170],seed[1004],seed[1844],seed[3402],seed[2841],seed[4046],seed[3289],seed[3729],seed[2037],seed[3691],seed[2845],seed[2663],seed[2321],seed[2302],seed[1135],seed[1694],seed[730],seed[3739],seed[3771],seed[2670],seed[838],seed[3598],seed[1229],seed[1820],seed[2716],seed[2272],seed[378],seed[1759],seed[3052],seed[1183],seed[444],seed[3411],seed[4002],seed[467],seed[3227],seed[3298],seed[1978],seed[3396],seed[2507],seed[1982],seed[2085],seed[53],seed[1012],seed[3629],seed[3882],seed[3190],seed[189],seed[974],seed[3476],seed[2766],seed[1778],seed[3672],seed[976],seed[2338],seed[1121],seed[4021],seed[3726],seed[1478],seed[3464],seed[1609],seed[2960],seed[3352],seed[1586],seed[222],seed[2634],seed[1380],seed[2121],seed[539],seed[3032],seed[3618],seed[2254],seed[940],seed[3589],seed[387],seed[2813],seed[283],seed[2363],seed[1994],seed[1508],seed[4069],seed[2392],seed[145],seed[3221],seed[2413],seed[3103],seed[3543],seed[1617],seed[1159],seed[1591],seed[704],seed[1811],seed[2750],seed[3948],seed[2978],seed[644],seed[1692],seed[2547],seed[3926],seed[2709],seed[989],seed[1990],seed[3850],seed[3255],seed[790],seed[2933],seed[3987],seed[758],seed[2370],seed[3340],seed[2452],seed[2045],seed[504],seed[2350],seed[715],seed[1944],seed[249],seed[2954],seed[3189],seed[3802],seed[2584],seed[3774],seed[3787],seed[3657],seed[1891],seed[1002],seed[1957],seed[3172],seed[2164],seed[182],seed[1096],seed[2444],seed[107],seed[137],seed[1866],seed[3886],seed[516],seed[3366],seed[3378],seed[3864],seed[2929],seed[1932],seed[2898],seed[2829],seed[1270],seed[1672],seed[2437],seed[847],seed[1986],seed[1246],seed[984],seed[1539],seed[1108],seed[2055],seed[3762],seed[900],seed[1429],seed[1136],seed[1663],seed[3659],seed[1186],seed[3855],seed[1298],seed[1205],seed[2014],seed[2504],seed[3307],seed[2857],seed[3846],seed[2245],seed[2724],seed[2990],seed[276],seed[762],seed[3082],seed[2679],seed[2449],seed[380],seed[2925],seed[3083],seed[776],seed[1352],seed[102],seed[3512],seed[239],seed[712],seed[1070],seed[3954],seed[1174],seed[470],seed[1378],seed[2889],seed[3747],seed[1860],seed[2764],seed[1633],seed[1871],seed[3563],seed[4066],seed[930],seed[313],seed[2489],seed[1921],seed[3213],seed[702],seed[477],seed[3637],seed[3317],seed[920],seed[1489],seed[148],seed[814],seed[752],seed[2318],seed[570],seed[75],seed[3471],seed[3090],seed[129],seed[1868],seed[3568],seed[2883],seed[2144],seed[118],seed[3288],seed[3640],seed[2839],seed[1943],seed[1143],seed[2969],seed[785],seed[2882],seed[933],seed[399],seed[1524],seed[2198],seed[2984],seed[3796],seed[3042],seed[2253],seed[3231],seed[3695],seed[511],seed[1430],seed[1885],seed[748],seed[2952],seed[2436],seed[1180],seed[156],seed[1559],seed[1410],seed[312],seed[464],seed[1592],seed[2049],seed[1936],seed[1032],seed[705],seed[1027],seed[3048],seed[14],seed[1590],seed[1796],seed[86],seed[3824],seed[1887],seed[3328],seed[416],seed[3047],seed[1545],seed[1114],seed[3239],seed[2975],seed[3452],seed[2789],seed[3521],seed[1749],seed[1991],seed[1359],seed[522],seed[1993],seed[3765],seed[1072],seed[2373],seed[1857],seed[1546],seed[1690],seed[1275],seed[2033],seed[1188],seed[2568],seed[1317],seed[2618],seed[2587],seed[2065],seed[3327],seed[1828],seed[1411],seed[913],seed[1766],seed[3952],seed[1001],seed[663],seed[476],seed[1630],seed[2794],seed[1181],seed[1449],seed[892],seed[978],seed[769],seed[2432],seed[3395],seed[3570],seed[1681],seed[3950],seed[1797],seed[1444],seed[3360],seed[1365],seed[496],seed[3781],seed[3078],seed[3522],seed[641],seed[319],seed[1098],seed[2887],seed[3144],seed[2869],seed[1752],seed[1798],seed[2548],seed[3936],seed[4082],seed[3021],seed[1819],seed[2273],seed[889],seed[1371],seed[544],seed[449],seed[2471],seed[3099],seed[2806],seed[446],seed[3119],seed[1011],seed[1669],seed[3062],seed[596],seed[1505],seed[383],seed[3313],seed[3012],seed[2953],seed[3937],seed[4016],seed[275],seed[3283],seed[3540],seed[1376],seed[3002],seed[1679],seed[2509],seed[166],seed[3000],seed[481],seed[729],seed[2745],seed[2596],seed[2374],seed[2554],seed[919],seed[607],seed[1392],seed[2067],seed[1462],seed[3872],seed[2078],seed[2397],seed[1735],seed[1916],seed[402],seed[471],seed[291],seed[2566],seed[1139],seed[165],seed[91],seed[2175],seed[135],seed[498],seed[1722],seed[3329],seed[1884],seed[1852],seed[2],seed[1008],seed[796],seed[1407],seed[4056],seed[1437],seed[1655],seed[3877],seed[1632],seed[1248],seed[3980],seed[3074],seed[2559],seed[2999],seed[1415],seed[3520],seed[524],seed[2830],seed[3400],seed[3755],seed[1848],seed[85],seed[1232],seed[3063],seed[1626],seed[2027],seed[1126],seed[202],seed[1329],seed[2783],seed[803],seed[508],seed[3995],seed[3219],seed[3717],seed[2398],seed[183],seed[263],seed[2438],seed[2294],seed[1439],seed[3694],seed[4012],seed[3176],seed[309],seed[2161],seed[49],seed[180],seed[1554],seed[458],seed[3891],seed[869],seed[2251],seed[1619],seed[3849],seed[3341],seed[3806],seed[1095],seed[1465],seed[1427],seed[927],seed[4087],seed[2997],seed[27],seed[3997],seed[1251],seed[285],seed[1925],seed[2900],seed[333],seed[3647],seed[343],seed[3264],seed[3656],seed[3704],seed[3690],seed[3139],seed[345],seed[2210],seed[1910],seed[2942],seed[2853],seed[1652],seed[2160],seed[3437],seed[3286],seed[2524],seed[2192],seed[868],seed[1556],seed[191],seed[3813],seed[32],seed[3611],seed[2972],seed[22],seed[4088],seed[622],seed[3669],seed[18],seed[909],seed[2316],seed[739],seed[3141],seed[649],seed[1241],seed[114],seed[1017],seed[2793],seed[891],seed[1306],seed[2415],seed[2215],seed[2620],seed[246],seed[3576],seed[104],seed[2785],seed[3727],seed[1227],seed[373],seed[3102],seed[2759],seed[1762],seed[3406],seed[2097],seed[1768],seed[3066],seed[3943],seed[1561],seed[422],seed[2863],seed[2303],seed[3990],seed[3157],seed[4052],seed[3949],seed[921],seed[3304],seed[2684],seed[4008],seed[1167],seed[2658],seed[844],seed[3868],seed[1544],seed[2178],seed[2649],seed[4011],seed[1036],seed[2629],seed[1280],seed[6],seed[1211],seed[3566],seed[3258],seed[3795],seed[2575],seed[1358],seed[2920],seed[3334],seed[4057],seed[451],seed[3092],seed[1051],seed[1454],seed[1000],seed[273],seed[723],seed[170],seed[3469],seed[1782],seed[3713],seed[2610],seed[3026],seed[1897],seed[2949],seed[1574],seed[3499],seed[751],seed[3638],seed[3243],seed[3041],seed[2693],seed[1696],seed[2203],seed[3785],seed[2106],seed[585],seed[119],seed[70],seed[2616],seed[228],seed[2451],seed[79],seed[355],seed[2747],seed[4079],seed[2331],seed[262],seed[975],seed[3683],seed[3551],seed[3034],seed[2054],seed[1510],seed[1644],seed[3965],seed[1418],seed[1423],seed[1729],seed[3971],seed[3662],seed[3851],seed[2001],seed[3594],seed[260],seed[794],seed[548],seed[3155],seed[1890],seed[3932],seed[1850],seed[1253],seed[1956],seed[216],seed[1784],seed[3423],seed[2878],seed[2569],seed[3491],seed[2797],seed[272],seed[1400],seed[1948],seed[1534],seed[2540],seed[763],seed[2112],seed[1294],seed[681],seed[3773],seed[3128],seed[2191],seed[3236],seed[3804],seed[2231],seed[3723],seed[3560],seed[232],seed[961],seed[2966],seed[3246],seed[3912],seed[2626],seed[3350],seed[2339],seed[1413],seed[3171],seed[1105],seed[2858],seed[303],seed[2140],seed[1573],seed[2523],seed[2276],seed[3974],seed[2199],seed[266],seed[822],seed[595],seed[1299],seed[1547],seed[3412],seed[3439],seed[1453],seed[115],seed[515],seed[861],seed[188],seed[634],seed[2760],seed[2039],seed[970],seed[92],seed[3652],seed[843],seed[297],seed[2156],seed[3985],seed[2943],seed[4076],seed[2257],seed[3351],seed[3383],seed[83],seed[1612],seed[2235],seed[3653],seed[3907],seed[3934],seed[3409],seed[3895],seed[3968],seed[2647],seed[3843],seed[7],seed[1041],seed[3096],seed[1414],seed[2940],seed[1014],seed[134],seed[2636],seed[4036],seed[998],seed[547],seed[4024],seed[1909],seed[96],seed[3956],seed[1970],seed[709],seed[2076],seed[1846],seed[2431],seed[3168],seed[2546],seed[2108],seed[980],seed[810],seed[2073],seed[2435],seed[2976],seed[3463],seed[3897],seed[1646],seed[485],seed[1757],seed[1841],seed[2007],seed[651],seed[1093],seed[1470],seed[1882],seed[2290],seed[125],seed[3725],seed[2287],seed[45],seed[3355],seed[35],seed[1417],seed[2383],seed[3832],seed[3532],seed[1110],seed[3530],seed[2499],seed[2248],seed[1285],seed[2711],seed[2926],seed[990],seed[1648],seed[2605],seed[3415],seed[2706],seed[3718],seed[384],seed[600],seed[3405],seed[3661],seed[2564],seed[307],seed[562],seed[2896],seed[2868],seed[2678],seed[2655],seed[825],seed[1397],seed[3731],seed[924],seed[2506],seed[999],seed[4034],seed[506],seed[3245],seed[1062],seed[1230],seed[1277],seed[2181],seed[2426],seed[1431],seed[3671],seed[1773],seed[4092],seed[1492],seed[4083],seed[459],seed[3805],seed[623],seed[4073],seed[2166],seed[167],seed[379],seed[828],seed[4078],seed[2744],seed[1319],seed[1747],seed[1926],seed[3545],seed[2704],seed[2577],seed[633],seed[362],seed[1588],seed[1101],seed[3468],seed[3507],seed[3558],seed[2842],seed[804],seed[944],seed[3754],seed[3248],seed[3478],seed[982],seed[3349],seed[1171],seed[3451],seed[3370],seed[201],seed[3195],seed[3104],seed[783],seed[826],seed[3939],seed[666],seed[1727],seed[679],seed[3076],seed[1687],seed[2638],seed[1447],seed[549],seed[1260],seed[3853],seed[2685],seed[1618],seed[3142],seed[1320],seed[3256],seed[1448],seed[2329],seed[3194]}; 
//        seed12 <= {seed[1889],seed[3760],seed[1435],seed[3054],seed[2990],seed[3895],seed[1623],seed[3431],seed[1622],seed[3944],seed[1128],seed[2206],seed[3167],seed[3857],seed[2912],seed[1789],seed[215],seed[691],seed[3978],seed[422],seed[957],seed[3940],seed[216],seed[1224],seed[3270],seed[2584],seed[696],seed[3293],seed[1049],seed[322],seed[3074],seed[1216],seed[3135],seed[386],seed[2041],seed[3005],seed[1720],seed[3133],seed[634],seed[1527],seed[2958],seed[2865],seed[2681],seed[966],seed[1436],seed[561],seed[876],seed[2549],seed[37],seed[1201],seed[485],seed[1582],seed[1169],seed[371],seed[301],seed[1648],seed[4002],seed[2062],seed[1108],seed[1865],seed[652],seed[1802],seed[3058],seed[272],seed[2233],seed[3197],seed[2184],seed[1199],seed[580],seed[1034],seed[3141],seed[158],seed[3151],seed[3343],seed[1876],seed[1331],seed[1411],seed[2575],seed[1072],seed[2477],seed[2017],seed[3313],seed[1430],seed[1237],seed[568],seed[1680],seed[2713],seed[3942],seed[1580],seed[665],seed[3998],seed[3236],seed[1280],seed[1801],seed[238],seed[2307],seed[3330],seed[2727],seed[1474],seed[1348],seed[2103],seed[2434],seed[3745],seed[3865],seed[3224],seed[826],seed[3291],seed[3811],seed[708],seed[2904],seed[821],seed[1235],seed[3856],seed[2698],seed[3644],seed[46],seed[2944],seed[1071],seed[4089],seed[2121],seed[3233],seed[2453],seed[3336],seed[3230],seed[2057],seed[1293],seed[3503],seed[2851],seed[1557],seed[401],seed[3273],seed[3264],seed[2197],seed[2693],seed[2910],seed[1499],seed[3189],seed[2678],seed[349],seed[1175],seed[1526],seed[3186],seed[3467],seed[2342],seed[1774],seed[436],seed[3366],seed[3108],seed[2075],seed[2525],seed[2625],seed[551],seed[3458],seed[3098],seed[1185],seed[1406],seed[1251],seed[3],seed[1725],seed[2523],seed[2791],seed[3826],seed[2080],seed[2319],seed[3539],seed[3154],seed[2170],seed[1603],seed[3408],seed[52],seed[1408],seed[2252],seed[889],seed[3164],seed[1518],seed[1891],seed[3551],seed[825],seed[2292],seed[520],seed[2399],seed[2038],seed[1536],seed[563],seed[2669],seed[1573],seed[2978],seed[1200],seed[1521],seed[1964],seed[3365],seed[3424],seed[2995],seed[3119],seed[3850],seed[21],seed[1745],seed[3791],seed[3731],seed[824],seed[2951],seed[3046],seed[2752],seed[4031],seed[521],seed[3742],seed[3908],seed[2943],seed[466],seed[2706],seed[3626],seed[412],seed[359],seed[4077],seed[2209],seed[90],seed[3001],seed[3957],seed[2949],seed[3461],seed[416],seed[2657],seed[1553],seed[290],seed[4039],seed[3795],seed[903],seed[441],seed[1697],seed[885],seed[3331],seed[3451],seed[2831],seed[3816],seed[1424],seed[455],seed[1578],seed[3846],seed[2249],seed[3335],seed[3262],seed[1286],seed[2253],seed[264],seed[2579],seed[2915],seed[3225],seed[3538],seed[2553],seed[1957],seed[3871],seed[60],seed[2665],seed[2235],seed[1857],seed[913],seed[1461],seed[3936],seed[2690],seed[3735],seed[3955],seed[1555],seed[3891],seed[2378],seed[103],seed[1595],seed[3641],seed[294],seed[526],seed[556],seed[2371],seed[2458],seed[3147],seed[2212],seed[245],seed[3199],seed[3642],seed[738],seed[1862],seed[904],seed[527],seed[1630],seed[1088],seed[1830],seed[2231],seed[312],seed[130],seed[395],seed[3607],seed[1223],seed[2430],seed[2815],seed[1144],seed[397],seed[3802],seed[1405],seed[1104],seed[1043],seed[3102],seed[2446],seed[2980],seed[1266],seed[3550],seed[3452],seed[2590],seed[848],seed[1998],seed[2333],seed[1395],seed[763],seed[1033],seed[1698],seed[2177],seed[2269],seed[410],seed[405],seed[2408],seed[3914],seed[2077],seed[3290],seed[2247],seed[2683],seed[4006],seed[263],seed[253],seed[1619],seed[3789],seed[658],seed[92],seed[1315],seed[757],seed[2884],seed[1272],seed[3268],seed[2410],seed[4082],seed[1150],seed[2945],seed[3276],seed[3041],seed[3966],seed[3591],seed[1139],seed[678],seed[991],seed[6],seed[2878],seed[1490],seed[4005],seed[995],seed[4020],seed[3967],seed[3980],seed[2830],seed[1911],seed[469],seed[2517],seed[1361],seed[1123],seed[1805],seed[2747],seed[2519],seed[3706],seed[667],seed[3127],seed[3298],seed[969],seed[2507],seed[370],seed[3606],seed[180],seed[609],seed[2159],seed[3462],seed[1611],seed[2028],seed[1415],seed[1892],seed[554],seed[1429],seed[666],seed[203],seed[3311],seed[4072],seed[91],seed[3316],seed[1218],seed[2597],seed[3919],seed[1585],seed[772],seed[1277],seed[3240],seed[3993],seed[1012],seed[2628],seed[2297],seed[127],seed[449],seed[3410],seed[472],seed[3786],seed[73],seed[417],seed[2711],seed[2930],seed[163],seed[1899],seed[3718],seed[1559],seed[2210],seed[3694],seed[1058],seed[2667],seed[2610],seed[2435],seed[3488],seed[484],seed[3161],seed[523],seed[2604],seed[3571],seed[3960],seed[2006],seed[854],seed[880],seed[1810],seed[1133],seed[3977],seed[2725],seed[599],seed[3125],seed[733],seed[140],seed[2736],seed[2056],seed[3035],seed[3471],seed[3509],seed[3725],seed[861],seed[289],seed[67],seed[3738],seed[3754],seed[3665],seed[1079],seed[1303],seed[2534],seed[898],seed[1860],seed[1078],seed[795],seed[1824],seed[2709],seed[4028],seed[126],seed[1843],seed[3817],seed[593],seed[4015],seed[2989],seed[850],seed[1628],seed[1528],seed[994],seed[1186],seed[2443],seed[2364],seed[2244],seed[4093],seed[1649],seed[2360],seed[2417],seed[1180],seed[3423],seed[2198],seed[2139],seed[11],seed[2708],seed[4085],seed[128],seed[2528],seed[1492],seed[3118],seed[3672],seed[3689],seed[549],seed[1929],seed[25],seed[1846],seed[2465],seed[1909],seed[2536],seed[618],seed[2354],seed[1346],seed[1096],seed[1325],seed[3324],seed[1294],seed[934],seed[204],seed[746],seed[2243],seed[1692],seed[2302],seed[1829],seed[1716],seed[74],seed[547],seed[1941],seed[3958],seed[145],seed[3381],seed[2228],seed[2048],seed[1335],seed[3649],seed[2167],seed[1242],seed[3755],seed[2343],seed[3003],seed[2758],seed[3299],seed[1020],seed[3409],seed[646],seed[1153],seed[2415],seed[1520],seed[2000],seed[1141],seed[3403],seed[1493],seed[85],seed[2969],seed[751],seed[985],seed[482],seed[305],seed[2270],seed[246],seed[1517],seed[2495],seed[684],seed[3188],seed[905],seed[2612],seed[356],seed[232],seed[2763],seed[468],seed[1779],seed[3620],seed[1589],seed[278],seed[2572],seed[1212],seed[4063],seed[3357],seed[835],seed[3628],seed[423],seed[3375],seed[3066],seed[3938],seed[4084],seed[1664],seed[2786],seed[2992],seed[3079],seed[3518],seed[3126],seed[1672],seed[3630],seed[2921],seed[1715],seed[641],seed[2405],seed[149],seed[1906],seed[4035],seed[3068],seed[2149],seed[595],seed[344],seed[1606],seed[292],seed[1481],seed[632],seed[3282],seed[1788],seed[3608],seed[2308],seed[793],seed[2923],seed[3781],seed[3541],seed[884],seed[3281],seed[2986],seed[681],seed[178],seed[385],seed[1885],seed[1130],seed[831],seed[2190],seed[40],seed[376],seed[133],seed[2412],seed[3807],seed[1285],seed[791],seed[2613],seed[1888],seed[1073],seed[2996],seed[944],seed[2794],seed[3542],seed[1412],seed[1060],seed[1665],seed[3612],seed[2275],seed[3679],seed[2259],seed[1143],seed[2451],seed[1349],seed[1304],seed[3768],seed[3269],seed[2288],seed[137],seed[1117],seed[1152],seed[516],seed[10],seed[2508],seed[3783],seed[2471],seed[328],seed[662],seed[2551],seed[2934],seed[2714],seed[1148],seed[3130],seed[1134],seed[3416],seed[3002],seed[477],seed[1399],seed[1605],seed[352],seed[3599],seed[788],seed[1763],seed[2619],seed[1712],seed[853],seed[1897],seed[3711],seed[870],seed[3156],seed[3563],seed[1506],seed[2592],seed[94],seed[2658],seed[3229],seed[2036],seed[2805],seed[3976],seed[142],seed[2386],seed[2457],seed[3194],seed[1807],seed[2656],seed[1693],seed[1917],seed[64],seed[2204],seed[1933],seed[743],seed[2039],seed[1197],seed[1268],seed[2699],seed[3825],seed[3379],seed[1247],seed[1145],seed[1271],seed[3413],seed[175],seed[220],seed[1083],seed[2445],seed[300],seed[132],seed[4062],seed[2882],seed[1187],seed[2467],seed[752],seed[1566],seed[940],seed[2183],seed[1390],seed[3097],seed[768],seed[562],seed[1529],seed[434],seed[2274],seed[1753],seed[62],seed[3279],seed[3842],seed[3243],seed[4040],seed[2131],seed[3866],seed[148],seed[3280],seed[1136],seed[2479],seed[956],seed[1717],seed[2670],seed[1916],seed[3176],seed[1702],seed[1507],seed[3064],seed[2854],seed[2751],seed[3110],seed[34],seed[697],seed[2723],seed[13],seed[2807],seed[3090],seed[465],seed[989],seed[3992],seed[1831],seed[3572],seed[1161],seed[1063],seed[4017],seed[1240],seed[3227],seed[2128],seed[1749],seed[3247],seed[1950],seed[2558],seed[888],seed[3000],seed[1439],seed[2700],seed[14],seed[2361],seed[3892],seed[1385],seed[3534],seed[2540],seed[3592],seed[2810],seed[2648],seed[1784],seed[2340],seed[2710],seed[2685],seed[740],seed[700],seed[3007],seed[571],seed[1082],seed[3870],seed[3323],seed[1051],seed[1598],seed[3426],seed[1848],seed[2491],seed[491],seed[2188],seed[637],seed[2724],seed[1524],seed[1669],seed[2223],seed[2050],seed[922],seed[4049],seed[2054],seed[297],seed[3882],seed[1711],seed[1444],seed[3078],seed[1227],seed[1983],seed[1232],seed[1539],seed[2439],seed[1639],seed[1990],seed[1821],seed[1914],seed[2022],seed[3739],seed[1509],seed[2127],seed[3748],seed[1599],seed[3277],seed[3080],seed[2178],seed[155],seed[2639],seed[1334],seed[1228],seed[2239],seed[2950],seed[3433],seed[3506],seed[1770],seed[2413],seed[3660],seed[654],seed[2688],seed[3931],seed[1955],seed[924],seed[820],seed[660],seed[3762],seed[1151],seed[3838],seed[2746],seed[3449],seed[2858],seed[2749],seed[2225],seed[4007],seed[1650],seed[467],seed[265],seed[3310],seed[2643],seed[965],seed[2011],seed[348],seed[3872],seed[745],seed[440],seed[3180],seed[2119],seed[3740],seed[3564],seed[3831],seed[343],seed[1569],seed[3082],seed[2144],seed[1695],seed[2448],seed[3019],seed[3470],seed[3637],seed[1744],seed[1627],seed[3474],seed[1996],seed[2913],seed[1262],seed[2888],seed[4019],seed[2599],seed[3445],seed[2407],seed[4034],seed[2087],seed[1236],seed[439],seed[2899],seed[3190],seed[1155],seed[2767],seed[2580],seed[2004],seed[2273],seed[3201],seed[3686],seed[2973],seed[3393],seed[570],seed[2015],seed[286],seed[584],seed[1596],seed[86],seed[2661],seed[1505],seed[3521],seed[711],seed[2102],seed[926],seed[3105],seed[972],seed[3034],seed[2256],seed[2304],seed[2433],seed[642],seed[3692],seed[45],seed[2023],seed[2692],seed[1985],seed[3766],seed[1905],seed[4080],seed[3528],seed[239],seed[2979],seed[4087],seed[1718],seed[1039],seed[3851],seed[2179],seed[494],seed[1401],seed[2780],seed[3926],seed[1122],seed[3884],seed[28],seed[897],seed[3578],seed[2920],seed[2005],seed[2328],seed[1340],seed[3049],seed[3537],seed[1626],seed[1095],seed[2608],seed[1781],seed[3193],seed[2109],seed[3719],seed[2030],seed[1523],seed[4073],seed[374],seed[535],seed[2373],seed[2897],seed[3833],seed[1026],seed[921],seed[2353],seed[1875],seed[3439],seed[3670],seed[3255],seed[2679],seed[935],seed[2018],seed[2376],seed[907],seed[3380],seed[2146],seed[1867],seed[2151],seed[1577],seed[3505],seed[2538],seed[3008],seed[110],seed[1488],seed[3805],seed[1545],seed[2444],seed[1561],seed[2120],seed[3210],seed[805],seed[3587],seed[3604],seed[3140],seed[2002],seed[727],seed[776],seed[2012],seed[2855],seed[1618],seed[3484],seed[1011],seed[3138],seed[1061],seed[1683],seed[2403],seed[3177],seed[1609],seed[2676],seed[1567],seed[1485],seed[497],seed[1041],seed[3069],seed[219],seed[1306],seed[3533],seed[1471],seed[3249],seed[2324],seed[458],seed[2492],seed[2694],seed[2089],seed[2909],seed[674],seed[167],seed[3038],seed[685],seed[3317],seed[933],seed[3026],seed[3989],seed[3737],seed[3651],seed[1883],seed[1930],seed[2890],seed[2073],seed[2626],seed[1312],seed[2422],seed[4004],seed[742],seed[3139],seed[760],seed[1548],seed[1787],seed[4044],seed[1313],seed[3655],seed[1961],seed[2152],seed[582],seed[3212],seed[3894],seed[3522],seed[895],seed[2115],seed[1057],seed[2021],seed[699],seed[1383],seed[1069],seed[2938],seed[1615],seed[3513],seed[2808],seed[669],seed[3111],seed[2594],seed[1901],seed[2],seed[1065],seed[2175],seed[3800],seed[3921],seed[1834],seed[3812],seed[1419],seed[2141],seed[592],seed[65],seed[2889],seed[2772],seed[2192],seed[3773],seed[3460],seed[1179],seed[2091],seed[1847],seed[2860],seed[3981],seed[2086],seed[1105],seed[29],seed[1602],seed[1106],seed[1691],seed[3367],seed[838],seed[1912],seed[2903],seed[27],seed[3621],seed[2827],seed[1341],seed[3114],seed[197],seed[3036],seed[460],seed[53],seed[533],seed[3923],seed[2722],seed[1017],seed[651],seed[2045],seed[3574],seed[3619],seed[3830],seed[3368],seed[1854],seed[2589],seed[3887],seed[3517],seed[522],seed[3597],seed[3933],seed[2695],seed[2562],seed[544],seed[256],seed[2305],seed[873],seed[1965],seed[1070],seed[1050],seed[1962],seed[2291],seed[2524],seed[2646],seed[2790],seed[2416],seed[190],seed[1005],seed[3319],seed[87],seed[3788],seed[1167],seed[815],seed[1554],seed[3158],seed[1677],seed[2237],seed[3615],seed[2485],seed[4067],seed[1337],seed[1953],seed[251],seed[1489],seed[2287],seed[2922],seed[3687],seed[529],seed[2759],seed[3875],seed[2497],seed[1927],seed[2985],seed[2647],seed[3456],seed[910],seed[2891],seed[3198],seed[892],seed[2964],seed[877],seed[3347],seed[2129],seed[2147],seed[2272],seed[2875],seed[3581],seed[1336],seed[611],seed[2455],seed[315],seed[2828],seed[1426],seed[2629],seed[2166],seed[3526],seed[2998],seed[1465],seed[61],seed[2777],seed[2283],seed[2560],seed[4074],seed[336],seed[1794],seed[1920],seed[2935],seed[3106],seed[1999],seed[3569],seed[2164],seed[3954],seed[1098],seed[3245],seed[1413],seed[2853],seed[369],seed[605],seed[2258],seed[3968],seed[1607],seed[1015],seed[1844],seed[1475],seed[1160],seed[3639],seed[2122],seed[2573],seed[41],seed[3478],seed[3720],seed[3053],seed[3905],seed[3318],seed[1305],seed[602],seed[2230],seed[3710],seed[655],seed[3787],seed[3705],seed[75],seed[616],seed[1328],seed[1783],seed[3836],seed[1101],seed[1456],seed[3314],seed[2196],seed[3004],seed[581],seed[3132],seed[3983],seed[3344],seed[2529],seed[2049],seed[229],seed[196],seed[3784],seed[420],seed[714],seed[836],seed[589],seed[1460],seed[2401],seed[3271],seed[66],seed[392],seed[3417],seed[799],seed[3384],seed[2662],seed[3415],seed[2263],seed[1402],seed[607],seed[247],seed[875],seed[2363],seed[1410],seed[2173],seed[623],seed[1149],seed[560],seed[47],seed[1102],seed[3822],seed[213],seed[1124],seed[2511],seed[3829],seed[3283],seed[3429],seed[1332],seed[649],seed[1931],seed[3045],seed[2927],seed[483],seed[2718],seed[868],seed[3308],seed[3399],seed[3839],seed[1678],seed[2214],seed[1719],seed[1841],seed[2883],seed[2817],seed[3202],seed[2555],seed[235],seed[2500],seed[172],seed[1881],seed[3238],seed[2279],seed[2541],seed[2505],seed[381],seed[1737],seed[3371],seed[3163],seed[1740],seed[3124],seed[2462],seed[950],seed[4051],seed[1296],seed[1183],seed[2241],seed[1252],seed[578],seed[2499],seed[4056],seed[1154],seed[273],seed[3912],seed[997],seed[150],seed[1202],seed[2917],seed[3434],seed[1255],seed[3083],seed[2084],seed[1441],seed[1035],seed[16],seed[983],seed[2418],seed[1519],seed[753],seed[1706],seed[1747],seed[368],seed[3761],seed[628],seed[2717],seed[871],seed[3500],seed[2929],seed[1945],seed[3267],seed[1701],seed[3376],seed[778],seed[722],seed[729],seed[2602],seed[4030],seed[3752],seed[3614],seed[594],seed[2886],seed[3671],seed[2901],seed[2208],seed[3169],seed[2754],seed[3350],seed[1068],seed[3730],seed[1882],seed[327],seed[2171],seed[785],seed[364],seed[20],seed[354],seed[4066],seed[1771],seed[2850],seed[3244],seed[3510],seed[144],seed[1376],seed[459],seed[3749],seed[451],seed[1416],seed[1014],seed[1915],seed[3094],seed[900],seed[786],seed[998],seed[100],seed[917],seed[1730],seed[3662],seed[1244],seed[2741],seed[2587],seed[489],seed[2372],seed[2298],seed[971],seed[4033],seed[2906],seed[928],seed[32],seed[2680],seed[1635],seed[3285],seed[230],seed[3585],seed[967],seed[2892],seed[902],seed[683],seed[307],seed[3855],seed[2156],seed[2470],seed[1168],seed[2282],seed[3454],seed[3172],seed[1006],seed[2172],seed[2516],seed[3516],seed[3485],seed[329],seed[1100],seed[908],seed[3329],seed[932],seed[2161],seed[139],seed[225],seed[4003],seed[1194],seed[3514],seed[1283],seed[2421],seed[3191],seed[2863],seed[1044],seed[1856],seed[1319],seed[3187],seed[4053],seed[1726],seed[1560],seed[310],seed[3647],seed[3373],seed[2094],seed[878],seed[1658],seed[1647],seed[3849],seed[182],seed[1594],seed[2406],seed[1620],seed[3322],seed[591],seed[1780],seed[3301],seed[3061],seed[704],seed[1025],seed[2357],seed[3498],seed[4050],seed[165],seed[3144],seed[1919],seed[4069],seed[268],seed[2707],seed[3043],seed[1980],seed[2644],seed[503],seed[1177],seed[3906],seed[1657],seed[3013],seed[3907],seed[3383],seed[2814],seed[226],seed[2955],seed[2180],seed[866],seed[2150],seed[942],seed[107],seed[1275],seed[3683],seed[2490],seed[2849],seed[2874],seed[1380],seed[915],seed[379],seed[1323],seed[2653],seed[1835],seed[2398],seed[961],seed[2603],seed[2240],seed[3530],seed[2303],seed[2033],seed[2003],seed[2313],seed[726],seed[2436],seed[3899],seed[2804],seed[3600],seed[576],seed[3214],seed[1450],seed[2203],seed[1687],seed[1090],seed[314],seed[2227],seed[2383],seed[83],seed[1353],seed[3820],seed[883],seed[2392],seed[1250],seed[3185],seed[2125],seed[1084],seed[2459],seed[3305],seed[3814],seed[1066],seed[3951],seed[1676],seed[672],seed[181],seed[698],seed[695],seed[1320],seed[3407],seed[3877],seed[3724],seed[2545],seed[1491],seed[3927],seed[3668],seed[1024],seed[1116],seed[3646],seed[2556],seed[511],seed[1081],seed[193],seed[138],seed[1111],seed[1616],seed[688],seed[1816],seed[3042],seed[2079],seed[1270],seed[2994],seed[2182],seed[1799],seed[1156],seed[2836],seed[3442],seed[2309],seed[759],seed[2335],seed[1951],seed[1479],seed[3237],seed[1302],seed[2800],seed[1734],seed[1356],seed[1671],seed[4047],seed[2290],seed[3695],seed[2673],seed[345],seed[63],seed[316],seed[1790],seed[1219],seed[1866],seed[3022],seed[920],seed[3027],seed[2503],seed[2099],seed[2654],seed[357],seed[1056],seed[3494],seed[762],seed[2637],seed[3726],seed[719],seed[214],seed[2677],seed[758],seed[2702],seed[3501],seed[3047],seed[1689],seed[3904],seed[1099],seed[2965],seed[1796],seed[1495],seed[2068],seed[3203],seed[4026],seed[1913],seed[1478],seed[2327],seed[3939],seed[3536],seed[1572],seed[1637],seed[1604],seed[811],seed[1556],seed[1873],seed[2696],seed[1688],seed[3263],seed[2916],seed[2861],seed[3840],seed[2911],seed[2475],seed[2820],seed[3174],seed[2729],seed[3780],seed[2472],seed[2261],seed[2163],seed[679],seed[1085],seed[1574],seed[2788],seed[1670],seed[1038],seed[1046],seed[675],seed[3885],seed[174],seed[510],seed[3828],seed[525],seed[3075],seed[2034],seed[781],seed[1022],seed[1516],seed[2530],seed[3702],seed[1995],seed[112],seed[1103],seed[2266],seed[114],seed[1992],seed[555],seed[2900],seed[2796],seed[1721],seed[960],seed[2756],seed[1273],seed[1817],seed[54],seed[3696],seed[3965],seed[2601],seed[566],seed[1513],seed[1284],seed[718],seed[1254],seed[702],seed[1295],seed[1203],seed[2104],seed[2348],seed[4012],seed[2130],seed[1003],seed[1125],seed[955],seed[3941],seed[2778],seed[3120],seed[3428],seed[1758],seed[2847],seed[689],seed[1469],seed[3232],seed[1984],seed[2533],seed[492],seed[1394],seed[1459],seed[2154],seed[2118],seed[2504],seed[3909],seed[659],seed[865],seed[744],seed[2844],seed[1354],seed[3974],seed[1409],seed[1925],seed[173],seed[993],seed[3476],seed[3611],seed[3018],seed[3845],seed[2420],seed[862],seed[919],seed[81],seed[3512],seed[2277],seed[1274],seed[1500],seed[1008],seed[2058],seed[860],seed[2856],seed[2873],seed[3582],seed[478],seed[1837],seed[129],seed[2264],seed[3101],seed[3360],seed[2789],seed[3395],seed[2926],seed[2521],seed[3136],seed[1142],seed[1887],seed[2512],seed[341],seed[2947],seed[3535],seed[1427],seed[1923],seed[2318],seed[1993],seed[1301],seed[2582],seed[3205],seed[1486],seed[2840],seed[3547],seed[2138],seed[2338],seed[3063],seed[51],seed[481],seed[1870],seed[2832],seed[3231],seed[3432],seed[1448],seed[1338],seed[687],seed[3767],seed[2060],seed[2400],seed[3020],seed[1926],seed[339],seed[4083],seed[3014],seed[3540],seed[822],seed[2771],seed[1575],seed[1979],seed[946],seed[2928],seed[1540],seed[3774],seed[1772],seed[2755],seed[3195],seed[2715],seed[400],seed[1404],seed[1714],seed[1989],seed[622],seed[2114],seed[2531],seed[2052],seed[453],seed[1037],seed[1166],seed[4029],seed[2143],seed[1674],seed[1681],seed[3048],seed[4070],seed[3583],seed[3307],seed[136],seed[1551],seed[1633],seed[378],seed[2966],seed[1751],seed[3779],seed[2522],seed[775],seed[1853],seed[627],seed[1795],seed[1653],seed[2332],seed[2195],seed[810],seed[615],seed[3995],seed[1047],seed[3584],seed[3295],seed[2255],seed[677],seed[3853],seed[3697],seed[4032],seed[38],seed[2615],seed[604],seed[1700],seed[2569],seed[3799],seed[2846],seed[2137],seed[1601],seed[1019],seed[620],seed[212],seed[210],seed[430],seed[121],seed[2914],seed[2098],seed[2552],seed[930],seed[280],seed[1898],seed[4048],seed[3459],seed[2450],seed[970],seed[108],seed[2869],seed[703],seed[2887],seed[1453],seed[2671],seed[3673],seed[3677],seed[3502],seed[2720],seed[3848],seed[518],seed[2359],seed[3753],seed[1221],seed[2801],seed[1207],seed[650],seed[1198],seed[818],seed[890],seed[118],seed[1921],seed[1769],seed[3148],seed[1852],seed[452],seed[1355],seed[2879],seed[3491],seed[1428],seed[2982],seed[3477],seed[1684],seed[160],seed[1591],seed[3093],seed[3463],seed[2924],seed[2339],seed[725],seed[1174],seed[2201],seed[2019],seed[1109],seed[852],seed[3032],seed[1859],seed[1818],seed[1703],seed[1510],seed[4013],seed[1278],seed[2806],seed[3159],seed[3055],seed[1241],seed[574],seed[285],seed[2781],seed[857],seed[279],seed[2219],seed[2257],seed[3804],seed[546],seed[539],seed[3192],seed[2750],seed[625],seed[3143],seed[1327],seed[415],seed[1009],seed[1625],seed[806],seed[1466],seed[1825],seed[4022],seed[3059],seed[567],seed[737],seed[626],seed[1590],seed[2107],seed[1127],seed[1632],seed[1982],seed[2775],seed[2007],seed[2390],seed[978],seed[323],seed[3092],seed[2894],seed[1994],seed[664],seed[3910],seed[3328],seed[3810],seed[2797],seed[84],seed[1021],seed[3402],seed[1359],seed[3801],seed[1248],seed[1414],seed[4046],seed[572],seed[864],seed[3364],seed[927],seed[2967],seed[3123],seed[2730],seed[3396],seed[396],seed[1075],seed[2194],seed[3566],seed[3699],seed[2682],seed[1814],seed[1205],seed[1791],seed[528],seed[2218],seed[3529],seed[260],seed[2632],seed[3028],seed[2948],seed[2145],seed[2812],seed[170],seed[3782],seed[1059],seed[1324],seed[3721],seed[2111],seed[1798],seed[2616],seed[1129],seed[701],seed[2396],seed[366],seed[1292],seed[977],seed[2083],seed[2042],seed[3287],seed[3504],seed[2867],seed[97],seed[2330],seed[2954],seed[1132],seed[3024],seed[3346],seed[3015],seed[2997],seed[1537],seed[1114],seed[2585],seed[918],seed[2380],seed[3631],seed[1903],seed[2454],seed[2460],seed[1864],seed[2704],seed[3656],seed[1833],seed[519],seed[2064],seed[517],seed[2893],seed[954],seed[1172],seed[3216],seed[1958],seed[332],seed[3349],seed[1112],seed[3924],seed[1115],seed[2957],seed[9],seed[2548],seed[1352],seed[346],seed[588],seed[3854],seed[244],seed[2488],seed[2550],seed[2798],seed[2618],seed[388],seed[179],seed[715],seed[373],seed[851],seed[3765],seed[779],seed[3095],seed[143],seed[2423],seed[721],seed[3837],seed[1329],seed[3552],seed[3261],seed[1952],seed[807],seed[1000],seed[3969],seed[1501],seed[2737],seed[1029],seed[77],seed[2481],seed[2323],seed[657],seed[1027],seed[2535],seed[1742],seed[33],seed[1815],seed[313],seed[1372],seed[2649],seed[4052],seed[1403],seed[887],seed[2331],seed[1288],seed[847],seed[2976],seed[406],seed[735],seed[1291],seed[456],seed[1690],seed[3217],seed[3573],seed[630],seed[269],seed[512],seed[2566],seed[2486],seed[1662],seed[2933],seed[3827],seed[3052],seed[2306],seed[4065],seed[2848],seed[4095],seed[2953],seed[3580],seed[1785],seed[30],seed[1624],seed[1544],seed[2666],seed[281],seed[2334],seed[3863],seed[199],seed[3181],seed[717],seed[1362],seed[1813],seed[3729],seed[841],seed[3627],seed[1682],seed[1384],seed[1822],seed[1535],seed[1257],seed[2296],seed[2735],seed[1258],seed[3691],seed[487],seed[790],seed[2972],seed[1502],seed[2547],seed[1373],seed[4009],seed[3722],seed[2742],seed[3325],seed[2819],seed[3684],seed[258],seed[564],seed[769],seed[43],seed[1126],seed[1016],seed[147],seed[1872],seed[19],seed[2782],seed[2356],seed[1565],seed[2464],seed[2761],seed[1253],seed[3128],seed[1608],seed[3618],seed[710],seed[3170],seed[2326],seed[2397],seed[3253],seed[1515],seed[3970],seed[2097],seed[3129],seed[794],seed[2440],seed[1457],seed[3497],seed[2384],seed[3440],seed[3254],seed[2574],seed[1863],seed[3868],seed[1991],seed[1970],seed[557],seed[1454],seed[2375],seed[540],seed[1612],seed[2478],seed[3411],seed[2543],seed[2442],seed[2870],seed[1091],seed[454],seed[3387],seed[3222],seed[3011],seed[1651],seed[1543],seed[3259],seed[168],seed[2857],seed[284],seed[2532],seed[1773],seed[3398],seed[2250],seed[186],seed[3418],seed[3985],seed[1724],seed[1417],seed[2135],seed[819],seed[464],seed[3678],seed[261],seed[399],seed[1775],seed[748],seed[1196],seed[2293],seed[1163],seed[3178],seed[241],seed[1443],seed[1811],seed[351],seed[404],seed[2544],seed[1778],seed[1571],seed[3950],seed[1287],seed[3242],seed[486],seed[96],seed[1260],seed[3659],seed[796],seed[2672],seed[2238],seed[3664],seed[1842],seed[4038],seed[1269],seed[3303],seed[2321],seed[78],seed[3115],seed[2085],seed[3155],seed[893],seed[48],seed[3466],seed[4042],seed[1425],seed[473],seed[2320],seed[1954],seed[712],seed[1389],seed[293],seed[3397],seed[1229],seed[3532],seed[2770],seed[899],seed[2093],seed[324],seed[2126],seed[541],seed[3545],seed[350],seed[986],seed[1878],seed[4008],seed[937],seed[2902],seed[923],seed[1377],seed[1256],seed[739],seed[3511],seed[1549],seed[783],seed[2301],seed[2743],seed[3771],seed[298],seed[2369],seed[1358],seed[3523],seed[3033],seed[499],seed[228],seed[3081],seed[1318],seed[1968],seed[2636],seed[3548],seed[1819],seed[1673],seed[1300],seed[680],seed[3629],seed[2381],seed[645],seed[3208],seed[2593],seed[3878],seed[1189],seed[1476],seed[1849],seed[1765],seed[1708],seed[131],seed[2035],seed[4037],seed[335],seed[3727],seed[3312],seed[610],seed[3815],seed[3386],seed[2082],seed[2826],seed[3076],seed[3337],seed[55],seed[2962],seed[803],seed[1587],seed[1210],seed[218],seed[2113],seed[3930],seed[2687],seed[1363],seed[2631],seed[2689],seed[1894],seed[1886],seed[1146],seed[377],seed[3309],seed[2181],seed[2868],seed[3601],seed[479],seed[509],seed[1048],seed[736],seed[3712],seed[1729],seed[3893],seed[988],seed[2939],seed[4018],seed[916],seed[2176],seed[3131],seed[2627],seed[2960],seed[1370],seed[488],seed[2617],seed[545],seed[2838],seed[1826],seed[3029],seed[614],seed[1614],seed[2026],seed[1741],seed[2200],seed[187],seed[1550],seed[827],seed[367],seed[3107],seed[1757],seed[1093],seed[3949],seed[200],seed[3874],seed[3218],seed[2385],seed[363],seed[421],seed[382],seed[3746],seed[2956],seed[2809],seed[3700],seed[387],seed[3602],seed[3353],seed[2222],seed[2701],seed[947],seed[3362],seed[1646],seed[2557],seed[3252],seed[2047],seed[2009],seed[3759],seed[217],seed[814],seed[2784],seed[2799],seed[3358],seed[2031],seed[1710],seed[2931],seed[437],seed[2216],seed[1067],seed[2919],seed[943],seed[797],seed[1137],seed[2576],seed[2732],seed[70],seed[3775],seed[360],seed[798],seed[912],seed[4010],seed[3717],seed[756],seed[3257],seed[3040],seed[3378],seed[471],seed[2733],seed[1343],seed[3603],seed[240],seed[3184],seed[2136],seed[4058],seed[2765],seed[3867],seed[843],seed[728],seed[2351],seed[1694],seed[3888],seed[361],seed[1445],seed[3421],seed[3847],seed[3294],seed[1282],seed[1823],seed[1713],seed[3085],seed[3616],seed[2651],seed[2981],seed[765],seed[1963],seed[2234],seed[3483],seed[3492],seed[1181],seed[2040],seed[693],seed[3663],seed[3226],seed[80],seed[3858],seed[2783],seed[1723],seed[1309],seed[2834],seed[288],seed[1446],seed[673],seed[692],seed[524],seed[1808],seed[31],seed[2907],seed[3685],seed[1939],seed[3643],seed[262],seed[1087],seed[1173],seed[1191],seed[390],seed[3579],seed[2088],seed[2559],seed[2571],seed[2368],seed[3559],seed[1666],seed[771],seed[159],seed[686],seed[3340],seed[2803],seed[237],seed[474],seed[375],seed[1298],seed[1345],seed[3165],seed[2586],seed[2614],seed[117],seed[640],seed[3852],seed[1977],seed[3961],seed[68],seed[2513],seed[1978],seed[2310],seed[3211],seed[1097],seed[3997],seed[1217],seed[1900],seed[3304],seed[1731],seed[3728],seed[3332],seed[1449],seed[3703],seed[2157],seed[3975],seed[2014],seed[855],seed[191],seed[2983],seed[538],seed[817],seed[925],seed[2456],seed[1761],seed[2076],seed[839],seed[408],seed[3900],seed[1877],seed[984],seed[2546],seed[317],seed[3590],seed[2463],seed[2630],seed[1514],seed[3793],seed[2987],seed[949],seed[3956],seed[1659],seed[2300],seed[1709],seed[3693],seed[4059],seed[3880],seed[3248],seed[590],seed[2224],seed[749],seed[2148],seed[2609],seed[1581],seed[1973],seed[3071],seed[2991],seed[254],seed[550],seed[2284],seed[1494],seed[3690],seed[3555],seed[3792],seed[151],seed[661],seed[7],seed[2065],seed[4079],seed[2285],seed[89],seed[2740],seed[1760],seed[2664],seed[3051],seed[1568],seed[2489],seed[980],seed[2668],seed[1231],seed[1064],seed[3100],seed[3420],seed[3701],seed[236],seed[2728],seed[3901],seed[1347],seed[829],seed[3708],seed[2936],seed[3681],seed[3050],seed[2016],seed[754],seed[3996],seed[1924],seed[1935],seed[2169],seed[2925],seed[2106],seed[1754],seed[1705],seed[36],seed[3286],seed[115],seed[3625],seed[2336],seed[3292],seed[583],seed[713],seed[3206],seed[504],seed[603],seed[1743],seed[2391],seed[716],seed[2074],seed[1052],seed[2642],seed[3289],seed[3932],seed[3757],seed[2349],seed[1470],seed[3577],seed[2606],seed[4060],seed[3351],seed[3635],seed[709],seed[906],seed[2051],seed[3864],seed[3750],seed[3088],seed[152],seed[413],seed[1832],seed[894],seed[93],seed[2294],seed[3982],seed[1746],seed[1442],seed[2165],seed[3457],seed[3117],seed[823],seed[495],seed[1290],seed[2611],seed[2946],seed[2063],seed[3374],seed[2311],seed[427],seed[4036],seed[2205],seed[3946],seed[833],seed[1080],seed[2101],seed[3918],seed[475],seed[3496],seed[3473],seed[2078],seed[3250],seed[2382],seed[2090],seed[1511],seed[3623],seed[2100],seed[1382],seed[1966],seed[1437],seed[3922],seed[221],seed[122],seed[3732],seed[207],seed[4025],seed[3468],seed[1643],seed[2600],seed[3438],seed[2236],seed[653],seed[2568],seed[629],seed[1645],seed[2501],seed[1592],seed[2426],seed[601],seed[2174],seed[3834],seed[3525],seed[3278],seed[2757],seed[1482],seed[4054],seed[2721],seed[1342],seed[2251],seed[3556],seed[1458],seed[515],seed[2289],seed[1316],seed[931],seed[3613],seed[4094],seed[1928],seed[3879],seed[362],seed[767],seed[962],seed[882],seed[3515],seed[979],seed[2242],seed[2968],seed[71],seed[1364],seed[3821],seed[222],seed[844],seed[2510],seed[619],seed[1264],seed[537],seed[1938],seed[1265],seed[3406],seed[3794],seed[3427],seed[867],seed[1388],seed[2880],seed[513],seed[1344],seed[101],seed[1699],seed[69],seed[3333],seed[1407],seed[3935],seed[2001],seed[891],seed[3808],seed[4],seed[3674],seed[1542],seed[1902],seed[3948],seed[3352],seed[548],seed[233],seed[1679],seed[3315],seed[2635],seed[1378],seed[1190],seed[1013],seed[2226],seed[1668],seed[2842],seed[2974],seed[3077],seed[3495],seed[3986],seed[419],seed[3334],seed[3401],seed[1367],seed[3044],seed[2248],seed[1946],seed[585],seed[231],seed[1934],seed[1001],seed[1944],seed[169],seed[3570],seed[1138],seed[4045],seed[3419],seed[3228],seed[176],seed[2476],seed[3796],seed[617],seed[2469],seed[4068],seed[1234],seed[2542],seed[257],seed[2494],seed[3898],seed[2108],seed[3756],seed[1634],seed[1121],seed[3297],seed[2142],seed[2813],seed[3062],seed[1861],seed[1238],seed[274],seed[1164],seed[2158],seed[879],seed[3806],seed[976],seed[3797],seed[2839],seed[125],seed[1040],seed[3321],seed[3785],seed[3012],seed[3251],seed[2341],seed[3508],seed[706],seed[3549],seed[2785],seed[2605],seed[3507],seed[1045],seed[1120],seed[1755],seed[1600],seed[3715],seed[22],seed[1431],seed[828],seed[3589],seed[945],seed[211],seed[2824],seed[1764],seed[1654],seed[3480],seed[1226],seed[2570],seed[383],seed[1800],seed[2387],seed[1895],seed[761],seed[613],seed[3113],seed[1546],seed[3593],seed[1766],seed[311],seed[3096],seed[2821],seed[1871],seed[15],seed[973],seed[340],seed[3447],seed[3223],seed[2337],seed[734],seed[1018],seed[104],seed[3680],seed[1728],seed[3650],seed[3609],seed[3889],seed[3070],seed[2908],seed[2134],seed[303],seed[2191],seed[1621],seed[308],seed[747],seed[177],seed[996],seed[4014],seed[3531],seed[2487],seed[1438],seed[3778],seed[1562],seed[3087],seed[1884],seed[1420],seed[3911],seed[44],seed[2262],seed[3487],seed[974],seed[3436],seed[975],seed[2554],seed[249],seed[3709],seed[201],seed[553],seed[2374],seed[141],seed[2872],seed[3881],seed[1113],seed[267],seed[389],seed[2211],seed[1947],seed[2823],seed[1062],seed[2719],seed[2971],seed[1597],seed[2008],seed[1496],seed[3675],seed[845],seed[1330],seed[2859],seed[188],seed[1195],seed[195],seed[2539],seed[2961],seed[2046],seed[2155],seed[2825],seed[3482],seed[801],seed[57],seed[2215],seed[2527],seed[670],seed[4075],seed[3073],seed[1777],seed[3122],seed[2703],seed[50],seed[444],seed[3037],seed[663],seed[2905],seed[3859],seed[705],seed[2932],seed[2186],seed[3657],seed[372],seed[302],seed[874],seed[3943],seed[1220],seed[2117],seed[2563],seed[2738],seed[1157],seed[959],seed[624],seed[1397],seed[1452],seed[438],seed[3764],seed[508],seed[1368],seed[3963],seed[3239],seed[2071],seed[3772],seed[3469],seed[2124],seed[447],seed[2059],seed[1748],seed[1004],seed[24],seed[3150],seed[3448],seed[1910],seed[3972],seed[4021],seed[326],seed[840],seed[3153],seed[2895],seed[1839],seed[3342],seed[536],seed[2013],seed[227],seed[1396],seed[333],seed[501],seed[1661],seed[1433],seed[1375],seed[774],seed[3869],seed[2473],seed[98],seed[2295],seed[1209],seed[2449],seed[2268],seed[3256],seed[1398],seed[3345],seed[3554],seed[3103],seed[3714],seed[3390],seed[2389],seed[2095],seed[981],seed[3913],seed[2774],seed[3450],seed[4078],seed[234],seed[1208],seed[896],seed[493],seed[787],seed[4023],seed[3776],seed[162],seed[1094],seed[3843],seed[4027],seed[2885],seed[3947],seed[2362],seed[939],seed[2634],seed[2760],seed[3196],seed[445],seed[2779],seed[3568],seed[3016],seed[2753],seed[3544],seed[1314],seed[470],seed[2140],seed[3372],seed[3617],seed[3744],seed[2940],seed[531],seed[3017],seed[3743],seed[3446],seed[506],seed[2822],seed[3741],seed[1140],seed[872],seed[1640],seed[2712],seed[171],seed[2344],seed[3896],seed[837],seed[2988],seed[586],seed[2975],seed[2480],seed[12],seed[1472],seed[3300],seed[3824],seed[2394],seed[1451],seed[2316],seed[476],seed[2072],seed[731],seed[2596],seed[2705],seed[1631],seed[3275],seed[1851],seed[4064],seed[2044],seed[2937],seed[1782],seed[2835],seed[2941],seed[1214],seed[543],seed[3654],seed[2502],seed[1736],seed[1279],seed[2744],seed[750],seed[3973],seed[682],seed[3798],seed[2187],seed[1162],seed[446],seed[3031],seed[3414],seed[2432],seed[276],seed[414],seed[59],seed[206],seed[3486],seed[2963],seed[1642],seed[2271],seed[1333],seed[1948],seed[26],seed[730],seed[1797],seed[304],seed[1440],seed[23],seed[3089],seed[1971],seed[3546],seed[3355],seed[259],seed[450],seed[1727],seed[1584],seed[2496],seed[2581],seed[1655],seed[1297],seed[1422],seed[2620],seed[909],seed[3272],seed[2025],seed[18],seed[2276],seed[2659],seed[35],seed[741],seed[2641],seed[2281],seed[2317],seed[2686],seed[3160],seed[2010],seed[3039],seed[3320],seed[1512],seed[498],seed[161],seed[135],seed[1213],seed[2918],seed[1768],seed[782],seed[3652],seed[500],seed[2787],seed[789],seed[1391],seed[1036],seed[418],seed[3475],seed[2474],seed[755],seed[1586],seed[849],seed[2280],seed[3713],seed[205],seed[1188],seed[3676],seed[812],seed[1667],seed[2466],seed[2484],seed[834],seed[3576],seed[1613],seed[3435],seed[2221],seed[2578],seed[2452],seed[1976],seed[3207],seed[2229],seed[1685],seed[3527],seed[255],seed[2246],seed[1263],seed[433],seed[1007],seed[156],seed[598],seed[3519],seed[1002],seed[3758],seed[1756],seed[2379],seed[119],seed[2768],seed[2818],seed[1969],seed[1350],seed[3220],seed[2776],seed[1733],seed[2871],seed[2583],seed[1360],seed[1534],seed[3937],seed[407],seed[3698],seed[3354],seed[1530],seed[2650],seed[2655],seed[2329],seed[2624],seed[3586],seed[1975],seed[4081],seed[2325],seed[3179],seed[1480],seed[1960],seed[530],seed[2793],seed[2053],seed[223],seed[2862],seed[1583],seed[384],seed[2567],seed[79],seed[2942],seed[2837],seed[596],seed[429],seed[3873],seed[355],seed[1357],seed[2069],seed[929],seed[2367],seed[3751],seed[3430],seed[111],seed[1868],seed[490],seed[542],seed[3520],seed[780],seed[558],seed[3453],seed[1423],seed[2621],seed[2055],seed[3288],seed[2260],seed[2745],seed[3183],seed[1786],seed[1563],seed[2267],seed[3175],seed[2366],seed[1178],seed[3084],seed[1176],seed[3091],seed[3567],seed[1735],seed[668],seed[3979],seed[1092],seed[3021],seed[3296],seed[3841],seed[2841],seed[2577],seed[3455],seed[1750],seed[275],seed[3769],seed[3356],seed[2388],seed[3803],seed[1076],seed[3723],seed[189],seed[3561],seed[2402],seed[1379],seed[1504],seed[2881],seed[1880],seed[3886],seed[3056],seed[2322],seed[1793],seed[2675],seed[3945],seed[1617],seed[2427],seed[3988],seed[1171],seed[3734],seed[3162],seed[309],seed[271],seed[1386],seed[3009],seed[2509],seed[3648],seed[1381],seed[2067],seed[3558],seed[2081],seed[1089],seed[1010],seed[3121],seed[3562],seed[277],seed[282],seed[773],seed[1317],seed[3030],seed[1579],seed[435],seed[1558],seed[1827],seed[116],seed[963],seed[443],seed[1547],seed[3575],seed[1365],seed[2811],seed[1576],seed[1387],seed[2358],seed[647],seed[2365],seed[2762],seed[941],seed[3633],seed[426],seed[804],seed[2565],seed[1467],seed[3987],seed[3359],seed[2189],seed[1552],seed[3876],seed[3274],seed[948],seed[331],seed[3400],seed[480],seed[3209],seed[120],seed[2734],seed[2286],seed[252],seed[3266],seed[1858],seed[1812],seed[1455],seed[2461],seed[2731],seed[1032],seed[154],seed[656],seed[39],seed[3200],seed[202],seed[987],seed[1762],seed[337],seed[3086],seed[2663],seed[2769],seed[1463],seed[194],seed[3543],seed[886],seed[707],seed[1806],seed[3704],seed[2561],seed[82],seed[1838],seed[2162],seed[1477],seed[411],seed[3391],seed[784],seed[3441],seed[1759],seed[2984],seed[1326],seed[2043],seed[1184],seed[1956],seed[1593],seed[3168],seed[1261],seed[911],seed[1042],seed[283],seed[3669],seed[1869],seed[321],seed[3023],seed[134],seed[4086],seed[724],seed[2483],seed[1588],seed[552],seed[1564],seed[358],seed[2876],seed[1525],seed[2185],seed[198],seed[951],seed[2748],seed[600],seed[992],seed[3844],seed[2520],seed[1828],seed[1222],seed[1722],seed[1652],seed[3658],seed[2112],seed[606],seed[3962],seed[3809],seed[569],seed[1988],seed[3394],seed[1322],seed[3991],seed[792],seed[3404],seed[2220],seed[3388],seed[3638],seed[266],seed[109],seed[2278],seed[2352],seed[635],seed[3006],seed[224],seed[1738],seed[2377],seed[1696],seed[3326],seed[1307],seed[2345],seed[502],seed[1893],seed[3109],seed[2447],seed[347],seed[2493],seed[3688],seed[3025],seed[1732],seed[3361],seed[1675],seed[2441],seed[1879],seed[1225],seed[587],seed[1054],seed[208],seed[105],seed[463],seed[3152],seed[1840],seed[2350],seed[1193],seed[2660],seed[1487],seed[1392],seed[3072],seed[1686],seed[1949],seed[2315],seed[1131],seed[106],seed[76],seed[3959],seed[1159],seed[325],seed[1211],seed[3443],seed[3425],seed[2977],seed[2370],seed[2414],seed[299],seed[1249],seed[1836],seed[802],seed[166],seed[2404],seed[1077],seed[2674],seed[1351],seed[4090],seed[639],seed[1767],seed[1192],seed[577],seed[1031],seed[3246],seed[442],seed[559],seed[2622],seed[1158],seed[3260],seed[846],seed[863],seed[2764],seed[2526],seed[3382],seed[800],seed[1170],seed[3284],seed[2697],seed[3104],seed[3137],seed[1922],seed[1739],seed[1610],seed[2845],seed[2970],seed[2037],seed[146],seed[968],seed[3917],seed[1369],seed[3883],seed[2096],seed[3707],seed[2061],seed[3265],seed[3925],seed[3984],seed[1028],seed[4000],seed[58],seed[2020],seed[964],seed[1],seed[2116],seed[319],seed[1165],seed[671],seed[2792],seed[49],seed[1147],seed[4016],seed[1497],seed[952],seed[2595],seed[2193],seed[3594],seed[3990],seed[2123],seed[2153],seed[3258],seed[3412],seed[1468],seed[1641],seed[1522],seed[2864],seed[2160],seed[3370],seed[1997],seed[1473],seed[3465],seed[859],seed[1937],seed[2691],seed[2070],seed[320],seed[2105],seed[2816],seed[124],seed[999],seed[72],seed[3823],seed[612],seed[2425],seed[3142],seed[380],seed[1023],seed[1803],seed[3481],seed[534],seed[365],seed[2029],seed[1447],seed[901],seed[3636],seed[1638],seed[2506],seed[1503],seed[914],seed[3971],seed[17],seed[1874],seed[631],seed[514],seed[3934],seed[690],seed[4055],seed[2202],seed[338],seed[1908],seed[1204],seed[2766],seed[573],seed[2355],seed[1118],seed[3770],seed[1629],seed[842],seed[2591],seed[608],seed[2419],seed[3437],seed[1371],seed[1418],seed[334],seed[3134],seed[1289],seed[2802],seed[644],seed[3112],seed[3479],seed[1393],seed[1644],seed[1896],seed[1245],seed[938],seed[1243],seed[1259],seed[764],seed[1972],seed[3790],seed[1532],seed[2232],seed[597],seed[3369],seed[3565],seed[1246],seed[393],seed[3338],seed[3595],seed[1321],seed[8],seed[496],seed[2092],seed[648],seed[3392],seed[1704],seed[3553],seed[808],seed[1374],seed[3489],seed[3166],seed[1400],seed[3661],seed[2999],seed[1776],seed[3302],seed[1940],seed[243],seed[2312],seed[2739],seed[1936],seed[2245],seed[2024],seed[398],seed[1918],seed[2393],seed[4057],seed[1311],seed[505],seed[1366],seed[123],seed[3099],seed[3813],seed[770],seed[2515],seed[1421],seed[816],seed[2428],seed[2429],seed[4011],seed[3835],seed[2623],seed[431],seed[3736],seed[242],seed[2346],seed[3405],seed[3377],seed[4076],seed[1432],seed[565],seed[3171],seed[2168],seed[1135],seed[425],seed[1974],seed[3929],seed[1986],seed[2110],seed[4001],seed[3624],seed[2716],seed[1086],seed[3903],seed[3385],seed[1981],seed[3348],seed[1792],seed[1959],seed[4061],seed[1541],seed[1904],seed[432],seed[1656],seed[296],seed[1498],seed[291],seed[507],seed[2199],seed[462],seed[3994],seed[3645],seed[4041],seed[3472],seed[2726],seed[1464],seed[1660],seed[402],seed[1890],seed[3234],seed[2437],seed[184],seed[4092],seed[3204],seed[3173],seed[2438],seed[3902],seed[953],seed[2795],seed[424],seed[295],seed[1119],seed[2898],seed[2431],seed[638],seed[1276],seed[394],seed[3596],seed[2314],seed[461],seed[3832],seed[1932],seed[3862],seed[1434],seed[3389],seed[3235],seed[2514],seed[3920],seed[2633],seed[403],seed[3640],seed[1230],seed[1281],seed[1570],seed[676],seed[2254],seed[3213],seed[1107],seed[3422],seed[2482],seed[2299],seed[3182],seed[982],seed[2066],seed[1310],seed[575],seed[3860],seed[99],seed[95],seed[766],seed[3666],seed[1339],seed[1707],seed[621],seed[990],seed[1206],seed[858],seed[3060],seed[4088],seed[1987],seed[830],seed[2607],seed[2027],seed[777],seed[157],seed[1804],seed[4091],seed[1943],seed[3861],seed[636],seed[2498],seed[1299],seed[2866],seed[448],seed[2133],seed[3818],seed[3634],seed[1053],seed[248],seed[643],seed[102],seed[2773],seed[3067],seed[330],seed[3747],seed[4024],seed[2217],seed[2959],seed[1855],seed[1845],seed[1308],seed[56],seed[3146],seed[3667],seed[3916],seed[1110],seed[2952],seed[3999],seed[3605],seed[1239],seed[2518],seed[4043],seed[1809],seed[3777],seed[869],seed[391],seed[3444],seed[723],seed[1233],seed[1752],seed[2833],seed[3964],seed[2213],seed[270],seed[1484],seed[2468],seed[3215],seed[633],seed[2265],seed[2411],seed[3341],seed[457],seed[318],seed[3897],seed[936],seed[2877],seed[1215],seed[113],seed[3588],seed[2409],seed[2032],seed[3327],seed[881],seed[88],seed[192],seed[2640],seed[809],seed[3219],seed[250],seed[409],seed[1483],seed[3363],seed[1967],seed[3010],seed[3610],seed[153],seed[3057],seed[3157],seed[0],seed[342],seed[1267],seed[4071],seed[1538],seed[2424],seed[1508],seed[183],seed[2537],seed[3763],seed[2645],seed[428],seed[2207],seed[2588],seed[732],seed[3632],seed[3953],seed[3560],seed[3682],seed[2829],seed[185],seed[2852],seed[579],seed[3499],seed[1663],seed[720],seed[2395],seed[353],seed[287],seed[532],seed[2993],seed[694],seed[1030],seed[2652],seed[3819],seed[42],seed[3464],seed[813],seed[1533],seed[856],seed[2347],seed[3149],seed[1636],seed[3890],seed[306],seed[1907],seed[3306],seed[2843],seed[958],seed[3557],seed[2598],seed[1820],seed[3241],seed[1182],seed[5],seed[3653],seed[2684],seed[3622],seed[3116],seed[3221],seed[2896],seed[164],seed[1074],seed[1462],seed[3952],seed[3524],seed[832],seed[3339],seed[3915],seed[3065],seed[3598],seed[1850],seed[209],seed[3493],seed[3733],seed[1531],seed[3490],seed[1942],seed[2564],seed[2132],seed[1055],seed[3145],seed[2638],seed[3716],seed[3928]};
//        seed13 <= {seed[2637],seed[694],seed[2721],seed[1265],seed[897],seed[3680],seed[2571],seed[1233],seed[866],seed[2447],seed[803],seed[536],seed[57],seed[827],seed[2742],seed[523],seed[305],seed[570],seed[1018],seed[33],seed[3448],seed[2408],seed[3419],seed[2792],seed[1566],seed[3413],seed[2068],seed[2167],seed[3122],seed[89],seed[1780],seed[1413],seed[3092],seed[858],seed[308],seed[2482],seed[2281],seed[2863],seed[251],seed[898],seed[855],seed[3575],seed[3080],seed[4023],seed[1322],seed[741],seed[149],seed[1258],seed[3555],seed[1677],seed[3383],seed[1578],seed[109],seed[3427],seed[1110],seed[2357],seed[239],seed[713],seed[3095],seed[309],seed[3628],seed[3664],seed[126],seed[379],seed[3140],seed[488],seed[1101],seed[3785],seed[3458],seed[3958],seed[3989],seed[2030],seed[3042],seed[103],seed[4020],seed[2595],seed[2188],seed[3604],seed[3607],seed[875],seed[2553],seed[1608],seed[260],seed[2183],seed[950],seed[1921],seed[359],seed[2265],seed[1557],seed[4039],seed[3154],seed[1231],seed[512],seed[2536],seed[147],seed[2170],seed[1889],seed[516],seed[2638],seed[915],seed[3250],seed[2052],seed[3356],seed[1073],seed[1562],seed[290],seed[3199],seed[2951],seed[2813],seed[2234],seed[1023],seed[3850],seed[3967],seed[3622],seed[3769],seed[697],seed[4043],seed[1296],seed[417],seed[1940],seed[792],seed[925],seed[3933],seed[1280],seed[2652],seed[276],seed[30],seed[2712],seed[2324],seed[3647],seed[3759],seed[3614],seed[1996],seed[3090],seed[1831],seed[2847],seed[1518],seed[1901],seed[2387],seed[2572],seed[3013],seed[2381],seed[2202],seed[2463],seed[157],seed[1136],seed[3948],seed[3873],seed[477],seed[2123],seed[232],seed[3313],seed[1631],seed[475],seed[1877],seed[1567],seed[1602],seed[1383],seed[2380],seed[220],seed[1686],seed[3502],seed[733],seed[1094],seed[2618],seed[2621],seed[3843],seed[775],seed[2740],seed[224],seed[2057],seed[3914],seed[375],seed[3959],seed[1708],seed[701],seed[911],seed[1180],seed[2133],seed[1038],seed[2418],seed[762],seed[1203],seed[1142],seed[2967],seed[254],seed[1432],seed[778],seed[1597],seed[568],seed[3477],seed[1282],seed[3827],seed[3161],seed[761],seed[184],seed[72],seed[228],seed[3976],seed[2020],seed[2707],seed[1556],seed[1834],seed[1174],seed[323],seed[98],seed[3182],seed[1781],seed[2877],seed[2431],seed[1320],seed[1793],seed[1181],seed[708],seed[1718],seed[1055],seed[3855],seed[2891],seed[3786],seed[441],seed[3815],seed[1267],seed[3936],seed[1473],seed[883],seed[2942],seed[2780],seed[4007],seed[1712],seed[3611],seed[1930],seed[2100],seed[3789],seed[3469],seed[1040],seed[2991],seed[3816],seed[2968],seed[1157],seed[1255],seed[979],seed[362],seed[110],seed[3739],seed[1010],seed[3303],seed[2625],seed[2474],seed[2770],seed[91],seed[2285],seed[3861],seed[3610],seed[3943],seed[1974],seed[3990],seed[1873],seed[661],seed[1008],seed[2500],seed[3652],seed[3937],seed[1962],seed[1495],seed[455],seed[1199],seed[2749],seed[2522],seed[2062],seed[1498],seed[3633],seed[1421],seed[2042],seed[2870],seed[2289],seed[2101],seed[3973],seed[3545],seed[798],seed[1293],seed[1559],seed[142],seed[1049],seed[2376],seed[404],seed[3314],seed[1388],seed[3075],seed[206],seed[1735],seed[3218],seed[3508],seed[3475],seed[2636],seed[3297],seed[526],seed[2475],seed[1170],seed[2941],seed[2731],seed[3594],seed[2643],seed[394],seed[1749],seed[696],seed[751],seed[3236],seed[3845],seed[2850],seed[2450],seed[4022],seed[2581],seed[1381],seed[1342],seed[2110],seed[175],seed[583],seed[808],seed[3134],seed[2327],seed[581],seed[3162],seed[2527],seed[3022],seed[6],seed[3331],seed[918],seed[3821],seed[1980],seed[3187],seed[2868],seed[386],seed[2141],seed[1493],seed[3328],seed[1818],seed[1364],seed[3893],seed[2488],seed[2258],seed[569],seed[1088],seed[2006],seed[2921],seed[3569],seed[557],seed[2095],seed[1738],seed[1347],seed[1403],seed[1987],seed[73],seed[1273],seed[3320],seed[2341],seed[2524],seed[3995],seed[3773],seed[69],seed[2270],seed[1279],seed[47],seed[2650],seed[90],seed[1451],seed[3077],seed[3979],seed[2689],seed[2913],seed[233],seed[2660],seed[182],seed[2144],seed[1066],seed[2119],seed[85],seed[92],seed[1097],seed[3412],seed[1439],seed[2084],seed[3846],seed[594],seed[3694],seed[108],seed[3919],seed[2980],seed[2125],seed[3315],seed[511],seed[1852],seed[352],seed[1392],seed[1540],seed[447],seed[3798],seed[3033],seed[1804],seed[2701],seed[61],seed[3782],seed[3517],seed[1574],seed[2292],seed[2129],seed[3145],seed[2746],seed[1747],seed[3925],seed[2287],seed[650],seed[1569],seed[2237],seed[2348],seed[373],seed[2074],seed[2458],seed[3568],seed[1946],seed[1515],seed[3209],seed[2692],seed[3668],seed[1299],seed[1437],seed[2817],seed[1806],seed[784],seed[498],seed[3757],seed[1648],seed[1820],seed[1630],seed[2412],seed[2319],seed[3868],seed[102],seed[508],seed[2768],seed[363],seed[3358],seed[3533],seed[912],seed[1799],seed[158],seed[2139],seed[3091],seed[3118],seed[873],seed[481],seed[29],seed[2539],seed[1212],seed[2986],seed[1918],seed[1898],seed[3345],seed[112],seed[3999],seed[2670],seed[948],seed[1828],seed[3335],seed[4008],seed[3509],seed[3360],seed[2704],seed[3440],seed[1645],seed[3120],seed[3932],seed[118],seed[757],seed[1797],seed[2711],seed[2104],seed[2714],seed[3210],seed[3205],seed[3025],seed[2912],seed[1007],seed[1655],seed[3691],seed[3586],seed[974],seed[3649],seed[1813],seed[544],seed[1976],seed[3423],seed[3188],seed[2212],seed[3211],seed[470],seed[3044],seed[1414],seed[3825],seed[947],seed[2346],seed[1458],seed[861],seed[1048],seed[3808],seed[2487],seed[848],seed[1098],seed[3130],seed[2051],seed[3975],seed[530],seed[1394],seed[2282],seed[3168],seed[1145],seed[3981],seed[2184],seed[2111],seed[395],seed[1395],seed[1721],seed[646],seed[2145],seed[351],seed[760],seed[2448],seed[2804],seed[3651],seed[237],seed[3201],seed[2113],seed[3666],seed[2869],seed[563],seed[2047],seed[3253],seed[288],seed[4001],seed[3867],seed[2254],seed[3641],seed[2858],seed[2932],seed[2723],seed[155],seed[2117],seed[41],seed[3831],seed[3325],seed[3333],seed[2922],seed[3219],seed[871],seed[1298],seed[1295],seed[2286],seed[1512],seed[2601],seed[3112],seed[83],seed[407],seed[1489],seed[2955],seed[1922],seed[944],seed[2541],seed[1288],seed[3105],seed[2271],seed[1917],seed[125],seed[1585],seed[3116],seed[2089],seed[1639],seed[2401],seed[3707],seed[2881],seed[926],seed[689],seed[3059],seed[436],seed[1925],seed[1244],seed[2058],seed[1990],seed[1125],seed[494],seed[2432],seed[4015],seed[1727],seed[3903],seed[1459],seed[1270],seed[3896],seed[2681],seed[2493],seed[1874],seed[1152],seed[657],seed[1189],seed[774],seed[221],seed[88],seed[3506],seed[3587],seed[200],seed[3483],seed[3035],seed[3371],seed[723],seed[3336],seed[1767],seed[905],seed[2366],seed[1651],seed[1341],seed[981],seed[2895],seed[1324],seed[687],seed[458],seed[3904],seed[2873],seed[1812],seed[3444],seed[3365],seed[921],seed[1571],seed[3052],seed[3408],seed[844],seed[319],seed[946],seed[3257],seed[3326],seed[1359],seed[1993],seed[2176],seed[2229],seed[2027],seed[3576],seed[1503],seed[2739],seed[1609],seed[2166],seed[3573],seed[2120],seed[2186],seed[261],seed[2717],seed[1740],seed[623],seed[1337],seed[2733],seed[339],seed[3504],seed[52],seed[2853],seed[3269],seed[1915],seed[3623],seed[3179],seed[1287],seed[4049],seed[3447],seed[3196],seed[549],seed[1286],seed[1128],seed[3086],seed[2426],seed[2677],seed[2501],seed[195],seed[2140],seed[3180],seed[1967],seed[1722],seed[1241],seed[879],seed[919],seed[1884],seed[1448],seed[1348],seed[3501],seed[138],seed[3947],seed[1516],seed[3629],seed[2776],seed[585],seed[3830],seed[695],seed[1688],seed[1961],seed[1469],seed[1294],seed[3701],seed[3688],seed[78],seed[3912],seed[137],seed[1719],seed[3512],seed[4014],seed[1254],seed[2800],seed[2886],seed[2259],seed[489],seed[2180],seed[2971],seed[2159],seed[2230],seed[1452],seed[3980],seed[2889],seed[3050],seed[3390],seed[2726],seed[66],seed[425],seed[133],seed[3388],seed[3391],seed[296],seed[3363],seed[3318],seed[727],seed[3164],seed[1785],seed[2112],seed[3375],seed[3535],seed[1202],seed[2196],seed[1616],seed[3171],seed[304],seed[1981],seed[3456],seed[3340],seed[439],seed[3415],seed[122],seed[3245],seed[1568],seed[3418],seed[360],seed[2065],seed[3730],seed[1118],seed[3395],seed[1752],seed[4086],seed[2861],seed[2149],seed[1166],seed[1120],seed[1851],seed[344],seed[592],seed[1580],seed[2339],seed[4012],seed[824],seed[3378],seed[144],seed[3791],seed[3818],seed[2856],seed[3264],seed[2702],seed[1237],seed[924],seed[2328],seed[1307],seed[2969],seed[1302],seed[2729],seed[53],seed[2246],seed[2538],seed[2419],seed[1988],seed[3767],seed[1809],seed[752],seed[3494],seed[1496],seed[411],seed[3076],seed[160],seed[1283],seed[2513],seed[940],seed[2175],seed[3765],seed[3716],seed[3638],seed[3267],seed[445],seed[95],seed[2083],seed[434],seed[448],seed[586],seed[3918],seed[1937],seed[1031],seed[759],seed[2152],seed[2477],seed[2273],seed[1576],seed[1702],seed[747],seed[2178],seed[719],seed[3811],seed[505],seed[665],seed[1973],seed[3372],seed[3015],seed[856],seed[1129],seed[484],seed[572],seed[2795],seed[3580],seed[2480],seed[2005],seed[3030],seed[2959],seed[2245],seed[1637],seed[259],seed[966],seed[3175],seed[1509],seed[2018],seed[2546],seed[3141],seed[982],seed[2761],seed[2405],seed[3554],seed[2478],seed[4072],seed[1099],seed[1113],seed[3528],seed[471],seed[1054],seed[2741],seed[3754],seed[2748],seed[1153],seed[3183],seed[1205],seed[3630],seed[3910],seed[2848],seed[870],seed[1778],seed[3747],seed[1084],seed[3496],seed[2250],seed[1319],seed[2266],seed[216],seed[1904],seed[1697],seed[2439],seed[3087],seed[2168],seed[1275],seed[2686],seed[4069],seed[1215],seed[217],seed[1433],seed[2845],seed[266],seed[653],seed[3146],seed[1707],seed[1162],seed[1005],seed[3834],seed[226],seed[630],seed[3058],seed[1528],seed[3272],seed[4077],seed[3480],seed[113],seed[2011],seed[2617],seed[3338],seed[3471],seed[4004],seed[1742],seed[3881],seed[189],seed[1179],seed[816],seed[1570],seed[1882],seed[4030],seed[3824],seed[1382],seed[3829],seed[2375],seed[1788],seed[1543],seed[3616],seed[1938],seed[614],seed[1680],seed[2841],seed[1713],seed[2197],seed[2545],seed[1530],seed[348],seed[4085],seed[2972],seed[2523],seed[989],seed[1687],seed[2658],seed[3278],seed[1832],seed[928],seed[3160],seed[3439],seed[26],seed[2404],seed[491],seed[3813],seed[1160],seed[3810],seed[1126],seed[4092],seed[4024],seed[1815],seed[2451],seed[185],seed[3273],seed[32],seed[2263],seed[2903],seed[3317],seed[2521],seed[401],seed[2803],seed[3312],seed[769],seed[2774],seed[2472],seed[4038],seed[3300],seed[2878],seed[1027],seed[4050],seed[1367],seed[2751],seed[3865],seed[190],seed[3887],seed[3069],seed[887],seed[3978],seed[3957],seed[952],seed[2081],seed[2876],seed[3485],seed[467],seed[3894],seed[954],seed[3064],seed[1720],seed[1075],seed[988],seed[515],seed[294],seed[2126],seed[63],seed[1711],seed[1067],seed[1971],seed[2824],seed[287],seed[1634],seed[1632],seed[1816],seed[3961],seed[616],seed[3492],seed[4010],seed[3942],seed[3531],seed[2198],seed[2283],seed[1551],seed[3909],seed[3429],seed[2135],seed[1186],seed[1600],seed[151],seed[2767],seed[1524],seed[3321],seed[3566],seed[1859],seed[3732],seed[3299],seed[909],seed[2840],seed[4047],seed[1610],seed[1964],seed[2732],seed[2516],seed[474],seed[524],seed[1091],seed[1340],seed[1256],seed[2703],seed[1150],seed[238],seed[793],seed[1879],seed[3343],seed[393],seed[114],seed[3561],seed[3579],seed[2849],seed[3449],seed[763],seed[1053],seed[4087],seed[1979],seed[148],seed[818],seed[3493],seed[2974],seed[1844],seed[1042],seed[613],seed[2148],seed[3734],seed[3750],seed[3593],seed[2954],seed[2326],seed[3702],seed[2651],seed[1857],seed[2679],seed[2910],seed[503],seed[256],seed[2044],seed[490],seed[2568],seed[100],seed[3800],seed[2189],seed[865],seed[3653],seed[183],seed[2818],seed[2136],seed[2305],seed[1044],seed[2407],seed[343],seed[1345],seed[50],seed[2243],seed[2709],seed[656],seed[3037],seed[2438],seed[336],seed[2543],seed[1374],seed[1969],seed[150],seed[1717],seed[3968],seed[3479],seed[746],seed[2783],seed[1855],seed[1537],seed[2471],seed[3753],seed[212],seed[850],seed[2037],seed[2008],seed[1449],seed[2616],seed[1856],seed[1491],seed[2436],seed[1285],seed[1513],seed[231],seed[755],seed[2984],seed[4091],seed[2570],seed[1725],seed[3807],seed[1849],seed[1590],seed[878],seed[2116],seed[3373],seed[3931],seed[1839],seed[1024],seed[3073],seed[3450],seed[2278],seed[2675],seed[671],seed[4074],seed[284],seed[1032],seed[3008],seed[3783],seed[2156],seed[1309],seed[560],seed[2316],seed[2187],seed[584],seed[1692],seed[3591],seed[198],seed[2288],seed[1396],seed[1850],seed[3403],seed[3525],seed[3115],seed[839],seed[2866],seed[428],seed[1245],seed[2452],seed[3156],seed[3268],seed[935],seed[19],seed[3900],seed[2384],seed[4002],seed[3776],seed[3292],seed[3377],seed[1490],seed[3930],seed[2620],seed[3128],seed[1953],seed[1910],seed[380],seed[3712],seed[2342],seed[1625],seed[3152],seed[649],seed[2907],seed[2276],seed[3203],seed[2661],seed[2730],seed[2309],seed[1483],seed[575],seed[3812],seed[2103],seed[3874],seed[3433],seed[501],seed[4036],seed[1249],seed[3571],seed[3287],seed[652],seed[76],seed[11],seed[2576],seed[3640],seed[3244],seed[1221],seed[1488],seed[1714],seed[3693],seed[2079],seed[662],seed[2077],seed[2397],seed[3157],seed[120],seed[2574],seed[2470],seed[4018],seed[84],seed[2777],seed[194],seed[1658],seed[1021],seed[1661],seed[1592],seed[1529],seed[3212],seed[885],seed[2865],seed[3728],seed[2540],seed[1045],seed[1681],seed[2585],seed[443],seed[4000],seed[2605],seed[2512],seed[3498],seed[3913],seed[209],seed[215],seed[2389],seed[3478],seed[2765],seed[922],seed[1734],seed[893],seed[163],seed[1071],seed[2495],seed[204],seed[459],seed[3537],seed[3663],seed[3240],seed[1028],seed[622],seed[3858],seed[3016],seed[3998],seed[3549],seed[2678],seed[1517],seed[2157],seed[4042],seed[881],seed[2925],seed[3070],seed[1754],seed[833],seed[1866],seed[3165],seed[749],seed[387],seed[3281],seed[642],seed[1497],seed[2952],seed[1876],seed[1875],seed[104],seed[3705],seed[250],seed[2093],seed[1934],seed[2799],seed[3768],seed[1078],seed[3167],seed[3715],seed[3801],seed[3627],seed[862],seed[3286],seed[2359],seed[1111],seed[1304],seed[4059],seed[1885],seed[1903],seed[3905],seed[107],seed[1694],seed[886],seed[3047],seed[2429],seed[976],seed[329],seed[2628],seed[2990],seed[3645],seed[680],seed[3302],seed[1746],seed[3686],seed[1363],seed[3305],seed[1741],seed[2199],seed[2299],seed[4057],seed[285],seed[242],seed[135],seed[2734],seed[2530],seed[1272],seed[2544],seed[2534],seed[2988],seed[3259],seed[1362],seed[1508],seed[1278],seed[2838],seed[1886],seed[3421],seed[1899],seed[1246],seed[1914],seed[1614],seed[2078],seed[2274],seed[2899],seed[12],seed[1739],seed[1002],seed[2242],seed[1191],seed[2191],seed[1243],seed[1116],seed[3396],seed[3382],seed[3],seed[2267],seed[1184],seed[2964],seed[229],seed[2607],seed[3949],seed[1108],seed[2713],seed[2331],seed[45],seed[2944],seed[3114],seed[3847],seed[998],seed[1888],seed[509],seed[571],seed[1554],seed[3578],seed[1823],seed[193],seed[1313],seed[1006],seed[1092],seed[235],seed[2473],seed[1536],seed[1138],seed[3654],seed[1555],seed[2798],seed[1628],seed[3956],seed[2094],seed[1505],seed[2115],seed[685],seed[2494],seed[2611],seed[202],seed[3915],seed[3232],seed[1761],seed[2771],seed[1972],seed[1195],seed[3696],seed[927],seed[3615],seed[2209],seed[655],seed[1955],seed[1081],seed[1864],seed[2306],seed[3697],seed[3362],seed[3608],seed[161],seed[2253],seed[3366],seed[1690],seed[2823],seed[2815],seed[754],seed[3417],seed[1957],seed[3039],seed[1247],seed[3227],seed[958],seed[1706],seed[3970],seed[3256],seed[543],seed[181],seed[3597],seed[1629],seed[2950],seed[3738],seed[620],seed[632],seed[410],seed[264],seed[3005],seed[821],seed[2039],seed[660],seed[2363],seed[500],seed[2185],seed[1626],seed[3246],seed[1748],seed[3006],seed[36],seed[553],seed[2846],seed[3529],seed[782],seed[2213],seed[1466],seed[2067],seed[3987],seed[1223],seed[96],seed[1709],seed[1698],seed[2926],seed[3177],seed[1956],seed[1867],seed[3637],seed[2710],seed[2313],seed[3584],seed[2232],seed[3612],seed[442],seed[3908],seed[369],seed[3662],seed[1519],seed[3119],seed[1950],seed[535],seed[2593],seed[3117],seed[1660],seed[3271],seed[2708],seed[3406],seed[1532],seed[3319],seed[1346],seed[1220],seed[3606],seed[2464],seed[2511],seed[3247],seed[74],seed[3195],seed[1595],seed[3658],seed[539],seed[1573],seed[3676],seed[403],seed[1970],seed[907],seed[3216],seed[2457],seed[366],seed[2296],seed[610],seed[809],seed[3027],seed[3735],seed[3720],seed[2097],seed[440],seed[3137],seed[3266],seed[1486],seed[1426],seed[2754],seed[328],seed[1482],seed[542],seed[1586],seed[1306],seed[1375],seed[1649],seed[3842],seed[2592],seed[580],seed[3283],seed[949],seed[303],seed[559],seed[3139],seed[2160],seed[3899],seed[2696],seed[2551],seed[178],seed[2904],seed[2936],seed[3742],seed[2307],seed[1531],seed[3285],seed[247],seed[2997],seed[2216],seed[3428],seed[293],seed[851],seed[3660],seed[2354],seed[2619],seed[1161],seed[3710],seed[2090],seed[3135],seed[3692],seed[3101],seed[838],seed[3397],seed[2608],seed[2982],seed[2021],seed[651],seed[3552],seed[2193],seed[628],seed[2315],seed[2531],seed[3648],seed[3558],seed[332],seed[771],seed[124],seed[270],seed[3675],seed[3851],seed[3771],seed[1881],seed[902],seed[1263],seed[2023],seed[546],seed[268],seed[2303],seed[2165],seed[2034],seed[3222],seed[207],seed[659],seed[277],seed[4065],seed[2872],seed[1615],seed[1906],seed[408],seed[2181],seed[3598],seed[1004],seed[1807],seed[3214],seed[146],seed[334],seed[959],seed[2888],seed[3011],seed[3826],seed[1544],seed[1526],seed[3426],seed[1100],seed[48],seed[1271],seed[2781],seed[418],seed[1774],seed[764],seed[188],seed[1646],seed[3174],seed[1253],seed[4066],seed[2340],seed[3736],seed[768],seed[3354],seed[2559],seed[2484],seed[2075],seed[2535],seed[1039],seed[548],seed[3169],seed[1082],seed[1547],seed[506],seed[4073],seed[3010],seed[3308],seed[492],seed[731],seed[1281],seed[1941],seed[337],seed[4089],seed[3155],seed[1926],seed[639],seed[22],seed[1389],seed[244],seed[996],seed[3526],seed[1998],seed[2409],seed[564],seed[1182],seed[132],seed[521],seed[2879],seed[307],seed[94],seed[1463],seed[3996],seed[888],seed[895],seed[1034],seed[3822],seed[3809],seed[3054],seed[116],seed[578],seed[3107],seed[4076],seed[579],seed[2312],seed[3237],seed[801],seed[396],seed[1290],seed[1035],seed[2355],seed[683],seed[1982],seed[1366],seed[811],seed[2134],seed[2802],seed[1456],seed[2343],seed[1619],seed[2885],seed[376],seed[3323],seed[1724],seed[3001],seed[2422],seed[2060],seed[1887],seed[3194],seed[1977],seed[2589],seed[111],seed[3066],seed[2639],seed[40],seed[3024],seed[3983],seed[3176],seed[3729],seed[3096],seed[3793],seed[3003],seed[1012],seed[2003],seed[1656],seed[34],seed[419],seed[2758],seed[1442],seed[2374],seed[1939],seed[882],seed[60],seed[3743],seed[2719],seed[2007],seed[1894],seed[3746],seed[3225],seed[599],seed[2421],seed[540],seed[27],seed[21],seed[3906],seed[3113],seed[3950],seed[829],seed[2855],seed[44],seed[278],seed[3724],seed[3596],seed[1783],seed[736],seed[3055],seed[2322],seed[514],seed[867],seed[1331],seed[3346],seed[3048],seed[1443],seed[1444],seed[169],seed[2364],seed[3466],seed[240],seed[3191],seed[3136],seed[1172],seed[3656],seed[1447],seed[1222],seed[3941],seed[1151],seed[3088],seed[3684],seed[2162],seed[3499],seed[814],seed[2820],seed[82],seed[799],seed[658],seed[3282],seed[3089],seed[1699],seed[2901],seed[2102],seed[1891],seed[2537],seed[997],seed[711],seed[758],seed[2793],seed[674],seed[370],seed[1905],seed[987],seed[1336],seed[1975],seed[218],seed[681],seed[4028],seed[3971],seed[1732],seed[3327],seed[1208],seed[438],seed[1323],seed[199],seed[1207],seed[3550],seed[2252],seed[3374],seed[720],seed[3885],seed[1214],seed[2498],seed[1771],seed[2467],seed[2843],seed[2909],seed[345],seed[2555],seed[3437],seed[1252],seed[3489],seed[3238],seed[2206],seed[4082],seed[1434],seed[4071],seed[3260],seed[537],seed[611],seed[1377],seed[3065],seed[1015],seed[2029],seed[2578],seed[1908],seed[3962],seed[3784],seed[4078],seed[3142],seed[2829],seed[1438],seed[3324],seed[2138],seed[706],seed[86],seed[2900],seed[3231],seed[1404],seed[1502],seed[702],seed[480],seed[1058],seed[2667],seed[3422],seed[2132],seed[1315],seed[3307],seed[1134],seed[3208],seed[1485],seed[1931],seed[971],seed[3491],seed[1504],seed[263],seed[1037],seed[2143],seed[2425],seed[1653],seed[1462],seed[2565],seed[3229],seed[3505],seed[3560],seed[3460],seed[1617],seed[325],seed[2688],seed[2588],seed[3543],seed[2241],seed[1096],seed[283],seed[2012],seed[728],seed[2264],seed[3452],seed[1830],seed[2054],seed[2778],seed[890],seed[2587],seed[2979],seed[3988],seed[51],seed[1117],seed[2836],seed[2646],seed[2987],seed[1399],seed[3602],seed[1301],seed[806],seed[3018],seed[2515],seed[3572],seed[740],seed[2382],seed[1772],seed[413],seed[3565],seed[3524],seed[364],seed[1511],seed[2875],seed[3751],seed[1932],seed[2594],seed[1453],seed[248],seed[615],seed[3657],seed[2529],seed[3060],seed[703],seed[357],seed[2573],seed[1072],seed[589],seed[1318],seed[174],seed[1642],seed[3643],seed[59],seed[3520],seed[3019],seed[1405],seed[2158],seed[469],seed[783],seed[933],seed[2017],seed[3454],seed[507],seed[551],seed[2221],seed[437],seed[555],seed[1520],seed[2000],seed[682],seed[1919],seed[3590],seed[2549],seed[2256],seed[2469],seed[2240],seed[2934],seed[3802],seed[2455],seed[4009],seed[1907],seed[2066],seed[4063],seed[291],seed[3953],seed[1095],seed[1327],seed[2064],seed[2235],seed[1836],seed[2417],seed[1123],seed[4090],seed[3002],seed[3848],seed[3974],seed[874],seed[286],seed[825],seed[3921],seed[1169],seed[3965],seed[1929],seed[2174],seed[2598],seed[3562],seed[2466],seed[2508],seed[734],seed[3511],seed[2718],seed[3659],seed[2687],seed[2414],seed[1696],seed[2356],seed[666],seed[3547],seed[2649],seed[3582],seed[1211],seed[637],seed[1542],seed[87],seed[3553],seed[3780],seed[518],seed[744],seed[1065],seed[2812],seed[1481],seed[127],seed[1158],seed[371],seed[3446],seed[1356],seed[3226],seed[1292],seed[1952],seed[3288],seed[392],seed[4095],seed[1057],seed[1784],seed[2153],seed[117],seed[3410],seed[3067],seed[300],seed[1026],seed[2244],seed[486],seed[1124],seed[2806],seed[1579],seed[1330],seed[3393],seed[3837],seed[3849],seed[612],seed[1693],seed[3760],seed[3669],seed[619],seed[4061],seed[1127],seed[1277],seed[1733],seed[2349],seed[2828],seed[3513],seed[820],seed[317],seed[576],seed[2410],seed[279],seed[1417],seed[3515],seed[2172],seed[1751],seed[3519],seed[341],seed[3166],seed[2514],seed[1763],seed[2070],seed[3839],seed[1352],seed[2373],seed[1043],seed[2350],seed[969],seed[208],seed[2706],seed[435],seed[3772],seed[3028],seed[3293],seed[2844],seed[3009],seed[2251],seed[698],seed[1627],seed[2906],seed[2599],seed[2096],seed[2329],seed[3451],seed[931],seed[16],seed[729],seed[673],seed[2561],seed[3261],seed[3945],seed[2837],seed[302],seed[957],seed[3880],seed[2519],seed[3476],seed[3852],seed[267],seed[2001],seed[1479],seed[1685],seed[213],seed[3193],seed[201],seed[3674],seed[1782],seed[1033],seed[2128],seed[1450],seed[3051],seed[1177],seed[2965],seed[3540],seed[4053],seed[1845],seed[1467],seed[1022],seed[454],seed[1548],seed[4068],seed[2632],seed[192],seed[2640],seed[1703],seed[3538],seed[795],seed[1052],seed[725],seed[3098],seed[1942],seed[18],seed[1726],seed[167],seed[2773],seed[942],seed[1470],seed[1471],seed[3392],seed[3523],seed[2489],seed[667],seed[2272],seed[910],seed[3764],seed[3626],seed[2736],seed[3123],seed[605],seed[1923],seed[2927],seed[863],seed[3866],seed[609],seed[3939],seed[2919],seed[269],seed[2295],seed[2669],seed[2291],seed[3275],seed[2962],seed[361],seed[3311],seed[1863],seed[1476],seed[2930],seed[2975],seed[624],seed[716],seed[1200],seed[2775],seed[776],seed[1606],seed[1549],seed[3559],seed[937],seed[2190],seed[2591],seed[3255],seed[3876],seed[787],seed[2961],seed[2600],seed[1912],seed[1730],seed[177],seed[2908],seed[1155],seed[627],seed[1076],seed[3097],seed[995],seed[3725],seed[1670],seed[1020],seed[281],seed[3796],seed[1563],seed[3964],seed[2437],seed[2918],seed[1840],seed[2610],seed[2154],seed[3721],seed[691],seed[1135],seed[1368],seed[608],seed[1829],seed[1985],seed[930],seed[2786],seed[1995],seed[3411],seed[1847],seed[2171],seed[714],seed[2108],seed[2393],seed[994],seed[1173],seed[934],seed[2635],seed[837],seed[153],seed[3886],seed[2146],seed[1525],seed[2105],seed[3871],seed[17],seed[3551],seed[289],seed[1872],seed[1425],seed[346],seed[4034],seed[3711],seed[1001],seed[3642],seed[3138],seed[1090],seed[1349],seed[2131],seed[1787],seed[1227],seed[826],seed[2],seed[2832],seed[4048],seed[3744],seed[3486],seed[3023],seed[3530],seed[3040],seed[450],seed[3034],seed[648],seed[4031],seed[1494],seed[2035],seed[4081],seed[3779],seed[1539],seed[3546],seed[943],seed[941],seed[128],seed[203],seed[2928],seed[3085],seed[1046],seed[872],seed[1700],seed[2896],seed[750],seed[3280],seed[25],seed[3698],seed[1657],seed[3198],seed[2043],seed[2092],seed[3963],seed[241],seed[2580],seed[2724],seed[415],seed[1361],seed[2998],seed[420],seed[960],seed[1080],seed[1623],seed[2978],seed[1933],seed[1289],seed[2905],seed[3589],seed[1800],seed[1764],seed[222],seed[565],seed[3761],seed[1682],seed[3683],seed[2563],seed[2280],seed[601],seed[2462],seed[3984],seed[186],seed[2575],seed[3386],seed[1947],seed[2835],seed[1596],seed[3790],seed[1750],seed[405],seed[721],seed[1613],seed[2630],seed[2400],seed[3817],seed[1790],seed[2890],seed[510],seed[381],seed[426],seed[1115],seed[3516],seed[1861],seed[2444],seed[3402],seed[678],seed[2238],seed[67],seed[3536],seed[1014],seed[1268],seed[3126],seed[2631],seed[3352],seed[3353],seed[1801],seed[2923],seed[173],seed[1047],seed[2325],seed[2031],seed[3869],seed[1621],seed[3057],seed[139],seed[39],seed[3290],seed[929],seed[1062],seed[1064],seed[2615],seed[3841],seed[2371],seed[2087],seed[903],seed[3111],seed[991],seed[2388],seed[3681],seed[2249],seed[37],seed[1167],seed[2973],seed[1593],seed[2490],seed[2048],seed[3541],seed[3709],seed[823],seed[301],seed[3084],seed[1779],seed[1729],seed[3892],seed[840],seed[1860],seed[0],seed[1365],seed[4021],seed[3110],seed[3158],seed[1089],seed[451],seed[1583],seed[457],seed[2874],seed[2779],seed[2173],seed[1997],seed[2526],seed[1197],seed[430],seed[1354],seed[65],seed[849],seed[3109],seed[1079],seed[3708],seed[3888],seed[93],seed[1016],seed[726],seed[1219],seed[1564],seed[1920],seed[2914],seed[3507],seed[965],seed[1407],seed[1674],seed[311],seed[2558],seed[1704],seed[2301],seed[2764],seed[115],seed[633],seed[2269],seed[3349],seed[4017],seed[1178],seed[1871],seed[1013],seed[1461],seed[1604],seed[3986],seed[3355],seed[2161],seed[3854],seed[3376],seed[3230],seed[3436],seed[236],seed[1063],seed[347],seed[917],seed[3603],seed[2690],seed[1140],seed[3459],seed[2468],seed[3241],seed[2496],seed[2685],seed[3472],seed[14],seed[1107],seed[868],seed[479],seed[3342],seed[2169],seed[1410],seed[906],seed[1441],seed[1499],seed[3197],seed[499],seed[1297],seed[28],seed[3689],seed[2333],seed[2697],seed[1343],seed[1011],seed[1507],seed[2217],seed[1880],seed[3254],seed[1500],seed[2377],seed[1652],seed[2107],seed[3178],seed[2787],seed[2204],seed[2528],seed[3733],seed[828],seed[2195],seed[3014],seed[1445],seed[1715],seed[900],seed[140],seed[1538],seed[2369],seed[3726],seed[2406],seed[2948],seed[3723],seed[1419],seed[3351],seed[836],seed[1546],seed[1335],seed[796],seed[834],seed[3857],seed[79],seed[2819],seed[449],seed[1984],seed[2737],seed[846],seed[1676],seed[3838],seed[669],seed[4005],seed[789],seed[901],seed[1777],seed[3994],seed[3737],seed[1131],seed[1429],seed[2399],seed[2441],seed[1316],seed[1753],seed[3079],seed[141],seed[1259],seed[1475],seed[522],seed[3316],seed[1406],seed[3190],seed[3542],seed[3289],seed[1662],seed[1228],seed[2810],seed[745],seed[832],seed[1059],seed[2569],seed[2360],seed[1669],seed[735],seed[629],seed[2378],seed[9],seed[590],seed[4019],seed[748],seed[1165],seed[3279],seed[3882],seed[2233],seed[3699],seed[3357],seed[3017],seed[3424],seed[2759],seed[62],seed[1112],seed[2634],seed[271],seed[3670],seed[1074],seed[772],seed[587],seed[2673],seed[2362],seed[986],seed[1792],seed[1386],seed[554],seed[797],seed[2834],seed[2791],seed[1185],seed[3159],seed[779],seed[472],seed[3147],seed[2808],seed[1594],seed[2228],seed[1892],seed[3094],seed[1527],seed[3510],seed[2150],seed[1262],seed[990],seed[1913],seed[3778],seed[2368],seed[1701],seed[3129],seed[4080],seed[4052],seed[1759],seed[282],seed[1371],seed[1843],seed[2036],seed[3220],seed[3124],seed[1510],seed[1959],seed[2454],seed[859],seed[3474],seed[1550],seed[2179],seed[1143],seed[800],seed[176],seed[2391],seed[1757],seed[3263],seed[1344],seed[647],seed[3398],seed[3379],seed[2231],seed[3213],seed[3527],seed[38],seed[2088],seed[4040],seed[1163],seed[1196],seed[2916],seed[2041],seed[321],seed[31],seed[2676],seed[2548],seed[3438],seed[2025],seed[399],seed[2788],seed[2811],seed[980],seed[1589],seed[2807],seed[465],seed[1853],seed[1902],seed[1019],seed[3488],seed[973],seed[3788],seed[3181],seed[1093],seed[179],seed[679],seed[2137],seed[1248],seed[3400],seed[3901],seed[327],seed[3056],seed[3004],seed[3977],seed[3775],seed[2365],seed[2668],seed[2109],seed[1858],seed[3667],seed[4093],seed[1821],seed[2069],seed[162],seed[2086],seed[2520],seed[493],seed[2337],seed[972],seed[654],seed[1665],seed[545],seed[664],seed[1620],seed[2983],seed[354],seed[595],seed[400],seed[1376],seed[805],seed[1384],seed[3291],seed[1171],seed[2935],seed[1387],seed[1314],seed[3934],seed[4079],seed[1762],seed[1041],seed[310],seed[1036],seed[1198],seed[3482],seed[1353],seed[984],seed[382],seed[223],seed[130],seed[3131],seed[3407],seed[780],seed[1009],seed[2633],seed[1003],seed[1415],seed[876],seed[342],seed[3828],seed[1737],seed[2411],seed[3405],seed[1083],seed[3370],seed[1402],seed[853],seed[1149],seed[2933],seed[2728],seed[444],seed[534],seed[1176],seed[2260],seed[3954],seed[738],seed[1795],seed[1427],seed[2506],seed[983],seed[358],seed[2782],seed[3186],seed[2533],seed[2827],seed[2222],seed[3441],seed[3875],seed[272],seed[3464],seed[1514],seed[1187],seed[3068],seed[3644],seed[2361],seed[978],seed[3548],seed[2999],seed[3745],seed[742],seed[923],seed[2814],seed[2497],seed[3920],seed[70],seed[2977],seed[1808],seed[2080],seed[2071],seed[743],seed[556],seed[3367],seed[2821],seed[4056],seed[2130],seed[1577],seed[2945],seed[1647],seed[626],seed[889],seed[3339],seed[2567],seed[81],seed[1264],seed[340],seed[1379],seed[2403],seed[1385],seed[3969],seed[3294],seed[1796],seed[2981],seed[2015],seed[280],seed[2725],seed[1664],seed[3153],seed[1261],seed[1949],seed[2210],seed[3856],seed[2700],seed[275],seed[3322],seed[955],seed[3242],seed[1408],seed[1776],seed[1400],seed[1260],seed[2435],seed[1989],seed[1416],seed[2398],seed[1390],seed[737],seed[2920],seed[1224],seed[2427],seed[262],seed[1393],seed[15],seed[2597],seed[2372],seed[2318],seed[3361],seed[2483],seed[1883],seed[1106],seed[1477],seed[2924],seed[3661],seed[1226],seed[2755],seed[421],seed[1728],seed[2353],seed[1193],seed[2279],seed[880],seed[412],seed[2525],seed[164],seed[3714],seed[2883],seed[1468],seed[1360],seed[1636],seed[1338],seed[3985],seed[2310],seed[456],seed[1339],seed[3381],seed[1274],seed[3359],seed[2182],seed[2939],seed[2902],seed[767],seed[54],seed[2680],seed[42],seed[602],seed[597],seed[3235],seed[2892],seed[1822],seed[1401],seed[2323],seed[717],seed[2367],seed[831],seed[2049],seed[2993],seed[577],seed[4083],seed[668],seed[3258],seed[625],seed[3401],seed[977],seed[318],seed[3570],seed[1744],seed[1909],seed[908],seed[2370],seed[3557],seed[365],seed[3104],seed[246],seed[462],seed[2949],seed[1317],seed[2666],seed[2004],seed[3063],seed[3026],seed[894],seed[2674],seed[2122],seed[292],seed[1936],seed[2698],seed[4027],seed[1060],seed[3585],seed[1201],seed[1994],seed[1087],seed[2050],seed[1325],seed[424],seed[3731],seed[3274],seed[1194],seed[4088],seed[3463],seed[24],seed[2826],seed[1133],seed[390],seed[2026],seed[2317],seed[3369],seed[1305],seed[2672],seed[2485],seed[2300],seed[2294],seed[2579],seed[985],seed[2505],seed[4045],seed[705],seed[2218],seed[3434],seed[3045],seed[2492],seed[2722],seed[3804],seed[1141],seed[4075],seed[1841],seed[3718],seed[3430],seed[1954],seed[3922],seed[1824],seed[2862],seed[2857],seed[1484],seed[2554],seed[1378],seed[2302],seed[2386],seed[1927],seed[1474],seed[3840],seed[429],seed[3583],seed[159],seed[1673],seed[2248],seed[3574],seed[1667],seed[3368],seed[1835],seed[1061],seed[1210],seed[3457],seed[1492],seed[2641],seed[3330],seed[4016],seed[3481],seed[1605],seed[2019],seed[672],seed[3740],seed[3248],seed[2583],seed[2352],seed[1944],seed[3631],seed[2024],seed[2655],seed[1587],seed[3567],seed[3020],seed[2642],seed[1572],seed[313],seed[1119],seed[4003],seed[830],seed[1945],seed[2268],seed[3619],seed[2032],seed[1575],seed[3394],seed[3766],seed[2192],seed[2211],seed[692],seed[2277],seed[2738],seed[3685],seed[1802],seed[106],seed[2970],seed[3618],seed[2992],seed[2214],seed[1817],seed[3532],seed[2604],seed[4067],seed[2164],seed[1916],seed[2629],seed[3836],seed[953],seed[1663],seed[97],seed[2790],seed[3748],seed[3207],seed[3897],seed[3252],seed[532],seed[3399],seed[1291],seed[3465],seed[932],seed[1350],seed[1644],seed[2127],seed[2224],seed[3284],seed[1321],seed[2747],seed[802],seed[566],seed[916],seed[2275],seed[432],seed[409],seed[1332],seed[1104],seed[1768],seed[1671],seed[3350],seed[2063],seed[2743],seed[2151],seed[904],seed[2720],seed[860],seed[80],seed[1535],seed[700],seed[3891],seed[338],seed[2963],seed[3484],seed[2860],seed[324],seed[1238],seed[813],seed[258],seed[1326],seed[55],seed[1758],seed[2772],seed[600],seed[3756],seed[3929],seed[3940],seed[274],seed[1069],seed[525],seed[2335],seed[3078],seed[473],seed[2091],seed[561],seed[3951],seed[1624],seed[3453],seed[3952],seed[1506],seed[2201],seed[1411],seed[1731],seed[538],seed[603],seed[71],seed[7],seed[2460],seed[2205],seed[3853],seed[1900],seed[2320],seed[773],seed[1188],seed[3133],seed[1983],seed[1423],seed[3173],seed[533],seed[676],seed[4041],seed[2753],seed[245],seed[168],seed[3081],seed[2830],seed[2960],seed[815],seed[2695],seed[1678],seed[2445],seed[3031],seed[520],seed[3072],seed[4064],seed[2582],seed[4037],seed[4055],seed[476],seed[2752],seed[1050],seed[3844],seed[896],seed[2624],seed[1598],seed[1239],seed[3883],seed[2550],seed[482],seed[2379],seed[297],seed[131],seed[2332],seed[2822],seed[2766],seed[641],seed[2219],seed[2756],seed[3955],seed[3102],seed[2566],seed[2220],seed[1372],seed[1056],seed[4046],seed[43],seed[3877],seed[1618],seed[964],seed[3895],seed[2385],seed[3409],seed[2225],seed[3083],seed[1370],seed[1465],seed[3923],seed[2613],seed[2509],seed[2098],seed[3234],seed[2453],seed[1560],seed[1541],seed[2654],seed[1965],seed[433],seed[383],seed[3521],seed[349],seed[463],seed[3306],seed[786],seed[3819],seed[3982],seed[2562],seed[1591],seed[4084],seed[3221],seed[2476],seed[3792],seed[3794],seed[2947],seed[1102],seed[1893],seed[1803],seed[2502],seed[961],seed[920],seed[2298],seed[1156],seed[3467],seed[2486],seed[2750],seed[2552],seed[2420],seed[372],seed[2801],seed[1068],seed[4054],seed[550],seed[631],seed[3495],seed[2481],seed[1232],seed[2659],seed[527],seed[3595],seed[2556],seed[3007],seed[2557],seed[3503],seed[2106],seed[3295],seed[1794],seed[3872],seed[2785],seed[3455],seed[2334],seed[2022],seed[2099],seed[3859],seed[2691],seed[3276],seed[3099],seed[3301],seed[2056],seed[2762],seed[3902],seed[13],seed[3993],seed[1743],seed[3599],seed[593],seed[842],seed[2082],seed[2255],seed[3935],seed[368],seed[1240],seed[753],seed[2479],seed[423],seed[1633],seed[693],seed[552],seed[817],seed[3556],seed[1229],seed[1723],seed[166],seed[2028],seed[1308],seed[2002],seed[1951],seed[790],seed[1948],seed[495],seed[2236],seed[3795],seed[333],seed[1357],seed[1168],seed[3564],seed[2745],seed[3490],seed[2590],seed[2118],seed[2059],seed[3189],seed[136],seed[1209],seed[2072],seed[2459],seed[99],seed[1148],seed[1588],seed[3884],seed[1789],seed[316],seed[388],seed[2794],seed[2033],seed[812],seed[1601],seed[822],seed[1561],seed[852],seed[2784],seed[219],seed[3749],seed[3462],seed[1668],seed[1454],seed[1234],seed[196],seed[3799],seed[732],seed[4011],seed[2396],seed[1355],seed[547],seed[3797],seed[1765],seed[519],seed[2851],seed[3106],seed[1077],seed[2648],seed[2958],seed[2989],seed[3144],seed[3924],seed[3082],seed[1825],seed[1827],seed[384],seed[2769],seed[191],seed[718],seed[2297],seed[962],seed[2416],seed[3577],seed[2816],seed[3832],seed[1760],seed[3148],seed[398],seed[1622],seed[3634],seed[2653],seed[2564],seed[992],seed[1978],seed[1643],seed[1218],seed[1358],seed[841],seed[1581],seed[3609],seed[1130],seed[496],seed[1373],seed[2428],seed[3310],seed[2744],seed[1869],seed[663],seed[3032],seed[1435],seed[2073],seed[3741],seed[3544],seed[1446],seed[640],seed[1862],seed[1786],seed[230],seed[618],seed[2392],seed[3385],seed[3200],seed[588],seed[3192],seed[1710],seed[3265],seed[2046],seed[2390],seed[677],seed[3108],seed[1798],seed[1154],seed[857],seed[847],seed[367],seed[330],seed[374],seed[3890],seed[210],seed[2940],seed[2684],seed[3991],seed[1329],seed[1159],seed[3814],seed[891],seed[1943],seed[2805],seed[1775],seed[3972],seed[3043],seed[1684],seed[406],seed[3348],seed[517],seed[312],seed[3687],seed[3468],seed[2560],seed[3960],seed[466],seed[3046],seed[574],seed[3755],seed[791],seed[1582],seed[3860],seed[2682],seed[1553],seed[2336],seed[1137],seed[1230],seed[2842],seed[2121],seed[617],seed[804],seed[2200],seed[1650],seed[715],seed[2657],seed[3497],seed[2893],seed[3296],seed[2596],seed[531],seed[2809],seed[143],seed[3170],seed[1928],seed[1654],seed[2124],seed[4070],seed[3927],seed[3805],seed[2957],seed[322],seed[1430],seed[356],seed[397],seed[119],seed[3600],seed[1000],seed[3944],seed[252],seed[1666],seed[788],seed[2434],seed[3431],seed[1896],seed[1086],seed[1250],seed[3387],seed[1791],seed[1303],seed[3781],seed[1584],seed[2344],seed[2953],seed[1412],seed[3601],seed[1819],seed[2946],seed[497],seed[3445],seed[1691],seed[1558],seed[2995],seed[3347],seed[607],seed[3966],seed[1689],seed[951],seed[558],seed[3143],seed[487],seed[4058],seed[1070],seed[2507],seed[2727],seed[154],seed[1351],seed[3916],seed[2938],seed[1312],seed[2395],seed[1999],seed[1183],seed[170],seed[56],seed[460],seed[75],seed[2456],seed[2311],seed[2010],seed[914],seed[10],seed[3997],seed[688],seed[845],seed[3000],seed[4013],seed[3695],seed[2215],seed[2290],seed[2994],seed[3341],seed[843],seed[1868],seed[3911],seed[3053],seed[709],seed[121],seed[2976],seed[3215],seed[295],seed[2239],seed[1085],seed[1029],seed[2898],seed[2662],seed[227],seed[645],seed[2894],seed[1679],seed[77],seed[1206],seed[1147],seed[591],seed[3270],seed[2911],seed[3416],seed[1276],seed[350],seed[2491],seed[2915],seed[739],seed[2884],seed[1814],seed[2014],seed[2937],seed[255],seed[1464],seed[3713],seed[2796],seed[2308],seed[2227],seed[385],seed[4035],seed[1310],seed[781],seed[1144],seed[1769],seed[2415],seed[567],seed[4094],seed[1640],seed[1960],seed[68],seed[2440],seed[1213],seed[187],seed[326],seed[869],seed[2917],seed[2394],seed[3404],seed[1409],seed[884],seed[2645],seed[502],seed[2797],seed[3870],seed[257],seed[3703],seed[3206],seed[2038],seed[1440],seed[452],seed[2735],seed[3679],seed[1242],seed[3514],seed[1192],seed[3803],seed[3621],seed[704],seed[1501],seed[1603],seed[562],seed[3889],seed[171],seed[1991],seed[3500],seed[2663],seed[3605],seed[3277],seed[2433],seed[234],seed[3617],seed[766],seed[4029],seed[2694],seed[298],seed[2155],seed[1146],seed[1534],seed[1391],seed[427],seed[3727],seed[596],seed[1225],seed[2226],seed[2897],seed[3364],seed[1755],seed[3635],seed[1472],seed[3719],seed[3636],seed[756],seed[2321],seed[1251],seed[2383],seed[3217],seed[1958],seed[1398],seed[2715],seed[1420],seed[3677],seed[2177],seed[1217],seed[1611],seed[3425],seed[3435],seed[416],seed[2586],seed[3700],seed[3938],seed[3823],seed[1457],seed[3149],seed[1328],seed[2358],seed[1257],seed[1051],seed[3150],seed[1565],seed[3062],seed[3470],seed[1109],seed[1418],seed[2402],seed[2854],seed[3121],seed[1216],seed[1736],seed[3334],seed[2055],seed[1612],seed[1854],seed[4006],seed[1],seed[3864],seed[2262],seed[3758],seed[864],seed[819],seed[3898],seed[1641],seed[4044],seed[2825],seed[2257],seed[2053],seed[2085],seed[2577],seed[1121],seed[1190],seed[1236],seed[1992],seed[320],seed[353],seed[2671],seed[635],seed[2223],seed[2430],seed[644],seed[3298],seed[3672],seed[3204],seed[3907],seed[152],seed[3038],seed[3673],seed[1030],seed[3613],seed[956],seed[1521],seed[2882],seed[3224],seed[3646],seed[2076],seed[2644],seed[2304],seed[165],seed[2996],seed[485],seed[3432],seed[1837],seed[1311],seed[2446],seed[724],seed[513],seed[1963],seed[3774],seed[2347],seed[3100],seed[1269],seed[1811],seed[3163],seed[3125],seed[2207],seed[180],seed[3682],seed[377],seed[1480],seed[105],seed[2833],seed[1460],seed[3946],seed[3127],seed[1204],seed[2504],seed[2852],seed[3690],seed[3380],seed[20],seed[3833],seed[3534],seed[1523],seed[3625],seed[5],seed[1164],seed[939],seed[1635],seed[2757],seed[3592],seed[2061],seed[1766],seed[1333],seed[3262],seed[2763],seed[1773],seed[3624],seed[3620],seed[2609],seed[1846],seed[2656],seed[638],seed[3563],seed[35],seed[3251],seed[730],seed[2443],seed[468],seed[634],seed[335],seed[3185],seed[315],seed[2532],seed[3172],seed[8],seed[3581],seed[2461],seed[3671],seed[2016],seed[145],seed[1745],seed[1132],seed[483],seed[606],seed[621],seed[1369],seed[464],seed[1695],seed[2518],seed[3632],seed[3704],seed[331],seed[835],seed[3442],seed[690],seed[765],seed[156],seed[391],seed[1838],seed[2956],seed[1848],seed[3806],seed[1533],seed[1675],seed[3588],seed[2716],seed[243],seed[2626],seed[49],seed[2867],seed[3243],seed[643],seed[3487],seed[686],seed[3706],seed[604],seed[2547],seed[3344],seed[402],seed[2943],seed[528],seed[3414],seed[4033],seed[2627],seed[253],seed[3863],seed[993],seed[3309],seed[1968],seed[134],seed[2985],seed[1284],seed[3539],seed[1175],seed[3021],seed[211],seed[1683],seed[355],seed[453],seed[4032],seed[1122],seed[794],seed[446],seed[3249],seed[2423],seed[699],seed[378],seed[3917],seed[3879],seed[810],seed[2664],seed[1017],seed[1870],seed[3835],seed[1716],seed[3443],seed[2647],seed[1545],seed[670],seed[1424],seed[2699],seed[129],seed[1599],seed[2147],seed[3132],seed[4026],seed[1607],seed[2194],seed[3678],seed[3461],seed[1431],seed[2351],seed[2864],seed[1428],seed[684],seed[1895],seed[2871],seed[3639],seed[3862],seed[478],seed[2831],seed[2208],seed[2887],seed[2693],seed[770],seed[899],seed[2839],seed[46],seed[2503],seed[1380],seed[2665],seed[1966],seed[1422],seed[2040],seed[1897],seed[2345],seed[2623],seed[3029],seed[1235],seed[2880],seed[197],seed[3420],seed[2510],seed[1924],seed[1266],seed[1025],seed[1842],seed[3992],seed[712],seed[2602],seed[2606],seed[1865],seed[2203],seed[892],seed[504],seed[1705],seed[877],seed[3228],seed[64],seed[2966],seed[3522],seed[2449],seed[2499],seed[573],seed[1935],seed[2603],seed[3202],seed[306],seed[461],seed[431],seed[722],seed[2705],seed[3820],seed[3928],seed[1890],seed[2612],seed[3787],seed[963],seed[3332],seed[3233],seed[1833],seed[2760],seed[1478],seed[1878],seed[3329],seed[1756],seed[2013],seed[214],seed[265],seed[975],seed[1139],seed[3103],seed[1455],seed[582],seed[807],seed[2789],seed[389],seed[3239],seed[3061],seed[4],seed[1300],seed[2330],seed[2424],seed[3041],seed[3337],seed[710],seed[2009],seed[777],seed[1810],seed[3752],seed[2465],seed[2931],seed[3049],seed[3071],seed[414],seed[2045],seed[2929],seed[785],seed[3650],seed[675],seed[2284],seed[101],seed[707],seed[1103],seed[2114],seed[3093],seed[1334],seed[3473],seed[23],seed[3184],seed[1397],seed[3389],seed[1672],seed[3926],seed[2142],seed[3722],seed[3036],seed[2584],seed[422],seed[3878],seed[205],seed[2413],seed[3384],seed[1770],seed[3770],seed[968],seed[3717],seed[249],seed[2859],seed[314],seed[1522],seed[2683],seed[529],seed[3151],seed[2261],seed[3665],seed[936],seed[854],seed[4025],seed[4051],seed[172],seed[1826],seed[1114],seed[970],seed[2517],seed[3074],seed[1638],seed[1986],seed[299],seed[3763],seed[1487],seed[1911],seed[2338],seed[4062],seed[3762],seed[1552],seed[273],seed[225],seed[1436],seed[938],seed[2442],seed[3223],seed[913],seed[2293],seed[2247],seed[2542],seed[999],seed[3304],seed[945],seed[3518],seed[1105],seed[2163],seed[2622],seed[1659],seed[3012],seed[598],seed[58],seed[2314],seed[636],seed[1805],seed[3655],seed[2614],seed[123],seed[3777],seed[541],seed[967],seed[4060]}; 
//        seed14 <= {seed[2718],seed[1655],seed[1349],seed[2651],seed[2271],seed[1920],seed[2133],seed[3033],seed[1147],seed[3493],seed[3143],seed[3813],seed[1282],seed[965],seed[2138],seed[3855],seed[1779],seed[2163],seed[3446],seed[1444],seed[109],seed[1414],seed[2943],seed[2341],seed[1598],seed[2033],seed[628],seed[2861],seed[1758],seed[3119],seed[2265],seed[2479],seed[3910],seed[271],seed[1139],seed[1006],seed[2361],seed[1930],seed[979],seed[91],seed[1843],seed[3617],seed[3190],seed[993],seed[2217],seed[2001],seed[3822],seed[873],seed[1510],seed[1924],seed[522],seed[612],seed[777],seed[1891],seed[757],seed[2219],seed[3352],seed[1218],seed[1348],seed[3199],seed[3260],seed[1576],seed[2537],seed[3373],seed[2956],seed[3018],seed[1462],seed[2522],seed[1820],seed[3148],seed[3688],seed[647],seed[3264],seed[2481],seed[1481],seed[365],seed[1938],seed[1752],seed[1411],seed[2004],seed[65],seed[2470],seed[4090],seed[3276],seed[501],seed[312],seed[3236],seed[939],seed[1571],seed[3080],seed[1525],seed[926],seed[3285],seed[1984],seed[764],seed[3680],seed[1328],seed[1251],seed[2516],seed[2258],seed[3667],seed[879],seed[872],seed[3379],seed[2659],seed[3126],seed[1508],seed[3381],seed[90],seed[1677],seed[2693],seed[3777],seed[7],seed[3610],seed[1181],seed[3637],seed[3189],seed[2740],seed[1352],seed[1237],seed[1198],seed[2419],seed[606],seed[14],seed[94],seed[1682],seed[2630],seed[2365],seed[1704],seed[2488],seed[1177],seed[2600],seed[2679],seed[1059],seed[914],seed[1472],seed[3521],seed[1199],seed[3991],seed[1337],seed[1153],seed[2552],seed[2994],seed[1267],seed[4016],seed[281],seed[3696],seed[2746],seed[421],seed[2327],seed[3536],seed[1997],seed[12],seed[3640],seed[2181],seed[3170],seed[294],seed[665],seed[1724],seed[517],seed[2476],seed[2967],seed[2503],seed[568],seed[1273],seed[2698],seed[3862],seed[3556],seed[2624],seed[1882],seed[1841],seed[592],seed[3642],seed[3205],seed[2287],seed[3280],seed[2373],seed[1538],seed[3097],seed[4051],seed[2836],seed[2834],seed[431],seed[2399],seed[3339],seed[2773],seed[1769],seed[2420],seed[3716],seed[1357],seed[2526],seed[3413],seed[1255],seed[384],seed[637],seed[713],seed[1464],seed[27],seed[3408],seed[135],seed[3055],seed[3215],seed[537],seed[2964],seed[3830],seed[2034],seed[383],seed[2066],seed[3449],seed[3477],seed[3098],seed[3090],seed[1520],seed[3155],seed[1903],seed[3824],seed[1913],seed[805],seed[1660],seed[656],seed[161],seed[3990],seed[661],seed[3041],seed[3917],seed[2543],seed[728],seed[1026],seed[2121],seed[1130],seed[3618],seed[3258],seed[2549],seed[268],seed[1917],seed[2412],seed[1263],seed[8],seed[802],seed[307],seed[2762],seed[1766],seed[3208],seed[2132],seed[3913],seed[1887],seed[3237],seed[1597],seed[604],seed[2865],seed[3432],seed[1961],seed[3766],seed[1505],seed[3218],seed[166],seed[120],seed[3300],seed[3374],seed[574],seed[538],seed[2665],seed[1032],seed[460],seed[3178],seed[2179],seed[2395],seed[1308],seed[652],seed[591],seed[2973],seed[617],seed[3593],seed[1848],seed[744],seed[3038],seed[3393],seed[704],seed[2821],seed[1854],seed[1523],seed[1201],seed[751],seed[1384],seed[2177],seed[3972],seed[2366],seed[1304],seed[1565],seed[3054],seed[2246],seed[413],seed[3816],seed[3590],seed[4026],seed[689],seed[2619],seed[1389],seed[500],seed[3282],seed[3130],seed[1594],seed[437],seed[916],seed[3011],seed[3865],seed[2403],seed[3516],seed[2962],seed[1974],seed[1128],seed[3158],seed[1784],seed[105],seed[1729],seed[3962],seed[1764],seed[3454],seed[2997],seed[1089],seed[1129],seed[718],seed[2433],seed[2013],seed[1585],seed[1686],seed[3946],seed[2256],seed[3444],seed[745],seed[2417],seed[29],seed[1725],seed[1787],seed[3140],seed[1007],seed[2368],seed[1477],seed[1539],seed[1794],seed[2996],seed[148],seed[3501],seed[2839],seed[3100],seed[2780],seed[1928],seed[3875],seed[2255],seed[2761],seed[2371],seed[302],seed[3682],seed[2618],seed[638],seed[1950],seed[723],seed[3572],seed[104],seed[4052],seed[1034],seed[385],seed[1061],seed[2335],seed[3240],seed[2176],seed[3228],seed[1722],seed[2095],seed[4003],seed[2782],seed[531],seed[1042],seed[3058],seed[3641],seed[2697],seed[2979],seed[382],seed[904],seed[84],seed[4070],seed[3294],seed[4009],seed[1781],seed[219],seed[3936],seed[2505],seed[2827],seed[284],seed[2666],seed[4005],seed[953],seed[3878],seed[2980],seed[1625],seed[3136],seed[1424],seed[511],seed[934],seed[3817],seed[3230],seed[1790],seed[836],seed[414],seed[1159],seed[3753],seed[3835],seed[3284],seed[1833],seed[2615],seed[3006],seed[3540],seed[1618],seed[3635],seed[3082],seed[3067],seed[1207],seed[1761],seed[3845],seed[1912],seed[1735],seed[3971],seed[1964],seed[1829],seed[3951],seed[1203],seed[3425],seed[110],seed[3307],seed[2143],seed[1617],seed[75],seed[2289],seed[3989],seed[3928],seed[2941],seed[454],seed[2506],seed[2447],seed[3330],seed[3639],seed[2146],seed[278],seed[308],seed[567],seed[554],seed[2750],seed[1688],seed[2885],seed[2038],seed[4014],seed[2749],seed[2947],seed[1856],seed[2915],seed[703],seed[1527],seed[3278],seed[2092],seed[1972],seed[3698],seed[3324],seed[1710],seed[2079],seed[425],seed[440],seed[206],seed[2111],seed[707],seed[4031],seed[2422],seed[1246],seed[3040],seed[3418],seed[1355],seed[3767],seed[851],seed[3726],seed[1036],seed[3973],seed[2064],seed[1316],seed[2999],seed[2873],seed[1786],seed[2633],seed[3654],seed[2021],seed[748],seed[597],seed[3009],seed[1692],seed[131],seed[3206],seed[2431],seed[1706],seed[2931],seed[528],seed[2350],seed[3792],seed[932],seed[1120],seed[1734],seed[898],seed[3160],seed[357],seed[2654],seed[903],seed[2290],seed[3281],seed[3725],seed[1543],seed[3029],seed[253],seed[3077],seed[1663],seed[2667],seed[2877],seed[215],seed[2923],seed[633],seed[3941],seed[2444],seed[927],seed[806],seed[1166],seed[1838],seed[601],seed[2691],seed[890],seed[2660],seed[2108],seed[2547],seed[2270],seed[3226],seed[1367],seed[185],seed[3219],seed[125],seed[60],seed[3386],seed[2778],seed[1522],seed[3524],seed[2957],seed[2316],seed[2074],seed[783],seed[840],seed[3378],seed[2484],seed[130],seed[1405],seed[2220],seed[1956],seed[349],seed[3626],seed[2497],seed[3305],seed[2105],seed[1172],seed[2715],seed[2527],seed[350],seed[2156],seed[328],seed[2449],seed[1380],seed[1802],seed[2360],seed[4019],seed[471],seed[406],seed[2813],seed[797],seed[2596],seed[158],seed[122],seed[3351],seed[1588],seed[1014],seed[180],seed[493],seed[1979],seed[3474],seed[4048],seed[313],seed[3153],seed[721],seed[3820],seed[2154],seed[96],seed[2791],seed[1043],seed[4006],seed[2427],seed[2211],seed[3052],seed[1814],seed[167],seed[1926],seed[648],seed[3580],seed[3288],seed[3037],seed[237],seed[3229],seed[2981],seed[3472],seed[2134],seed[2717],seed[121],seed[2195],seed[2560],seed[321],seed[3814],seed[182],seed[2758],seed[3883],seed[509],seed[2644],seed[2607],seed[2169],seed[3560],seed[1876],seed[20],seed[404],seed[828],seed[945],seed[174],seed[2508],seed[147],seed[825],seed[2533],seed[2261],seed[1792],seed[2765],seed[3597],seed[544],seed[1503],seed[1236],seed[2755],seed[543],seed[3712],seed[99],seed[3473],seed[1487],seed[3988],seed[1134],seed[2763],seed[1416],seed[3577],seed[4000],seed[1229],seed[552],seed[3721],seed[1743],seed[3089],seed[2187],seed[1087],seed[1124],seed[2523],seed[2472],seed[2022],seed[286],seed[98],seed[4035],seed[1874],seed[1708],seed[463],seed[2230],seed[176],seed[1002],seed[3411],seed[919],seed[2656],seed[822],seed[583],seed[782],seed[2393],seed[1277],seed[790],seed[1265],seed[3396],seed[2262],seed[881],seed[2223],seed[3749],seed[3841],seed[1826],seed[3387],seed[3921],seed[4037],seed[2385],seed[2392],seed[3670],seed[632],seed[3863],seed[513],seed[1537],seed[3484],seed[2482],seed[2952],seed[3558],seed[395],seed[1817],seed[1458],seed[423],seed[1433],seed[2315],seed[870],seed[126],seed[1687],seed[2298],seed[2905],seed[5],seed[1716],seed[2291],seed[3608],seed[3275],seed[1528],seed[2390],seed[3860],seed[265],seed[1593],seed[1944],seed[0],seed[2858],seed[1546],seed[288],seed[2308],seed[1100],seed[181],seed[1855],seed[3856],seed[1497],seed[2218],seed[3809],seed[3162],seed[2535],seed[2018],seed[1209],seed[2669],seed[407],seed[2539],seed[3684],seed[3853],seed[2306],seed[157],seed[1023],seed[1774],seed[1737],seed[3554],seed[856],seed[2463],seed[1090],seed[716],seed[2672],seed[1985],seed[1257],seed[3195],seed[3507],seed[3061],seed[3899],seed[2436],seed[1581],seed[3919],seed[2362],seed[3397],seed[2090],seed[2297],seed[3960],seed[1064],seed[1278],seed[2907],seed[2948],seed[3429],seed[3065],seed[3615],seed[2023],seed[2515],seed[3581],seed[2151],seed[175],seed[2448],seed[2793],seed[3812],seed[410],seed[2029],seed[3401],seed[3837],seed[762],seed[3606],seed[2716],seed[4057],seed[1286],seed[2052],seed[959],seed[3966],seed[603],seed[2728],seed[3548],seed[848],seed[865],seed[1048],seed[621],seed[277],seed[3768],seed[2859],seed[3594],seed[2234],seed[459],seed[2369],seed[2601],seed[3481],seed[3075],seed[640],seed[759],seed[332],seed[4013],seed[3673],seed[690],seed[4010],seed[3685],seed[82],seed[149],seed[1154],seed[1919],seed[2880],seed[3326],seed[267],seed[2807],seed[2326],seed[1501],seed[1805],seed[3629],seed[774],seed[4032],seed[521],seed[1270],seed[2511],seed[4073],seed[2178],seed[272],seed[818],seed[3166],seed[1951],seed[1310],seed[4007],seed[3665],seed[3415],seed[3889],seed[3131],seed[4002],seed[247],seed[2490],seed[3675],seed[455],seed[838],seed[3069],seed[949],seed[2838],seed[2707],seed[1183],seed[364],seed[3949],seed[2845],seed[3539],seed[3464],seed[2816],seed[3471],seed[1850],seed[2115],seed[264],seed[2574],seed[1696],seed[3181],seed[3430],seed[129],seed[4047],seed[3791],seed[666],seed[2123],seed[244],seed[3801],seed[670],seed[920],seed[1858],seed[1999],seed[1504],seed[1359],seed[1379],seed[2814],seed[2922],seed[1863],seed[2673],seed[3914],seed[266],seed[2280],seed[2235],seed[3360],seed[3727],seed[2440],seed[3839],seed[3492],seed[389],seed[1131],seed[2823],seed[518],seed[2453],seed[4075],seed[3745],seed[2008],seed[758],seed[2507],seed[361],seed[1605],seed[1676],seed[896],seed[588],seed[112],seed[2128],seed[2810],seed[2846],seed[3690],seed[34],seed[1822],seed[1506],seed[1670],seed[3840],seed[1055],seed[3161],seed[143],seed[3355],seed[1008],seed[3515],seed[1816],seed[3699],seed[33],seed[3347],seed[3505],seed[171],seed[231],seed[859],seed[2592],seed[1895],seed[2971],seed[3269],seed[2863],seed[3296],seed[1419],seed[769],seed[1213],seed[1327],seed[2227],seed[4017],seed[3409],seed[1610],seed[3895],seed[1775],seed[846],seed[2048],seed[3013],seed[2245],seed[676],seed[664],seed[2175],seed[2257],seed[3705],seed[2955],seed[3405],seed[426],seed[1275],seed[3969],seed[2379],seed[1215],seed[709],seed[381],seed[1493],seed[1910],seed[651],seed[2870],seed[275],seed[3701],seed[1170],seed[2414],seed[2556],seed[453],seed[3672],seed[529],seed[964],seed[204],seed[2058],seed[2895],seed[3894],seed[352],seed[1496],seed[2323],seed[2803],seed[784],seed[1550],seed[3297],seed[114],seed[826],seed[639],seed[921],seed[69],seed[1434],seed[1473],seed[3335],seed[3873],seed[1762],seed[2231],seed[1853],seed[2978],seed[1544],seed[2963],seed[3785],seed[2078],seed[1322],seed[3761],seed[297],seed[2321],seed[733],seed[958],seed[4067],seed[771],seed[2221],seed[1827],seed[2239],seed[2016],seed[3354],seed[3589],seed[1712],seed[3116],seed[1992],seed[2404],seed[2467],seed[1070],seed[3030],seed[3486],seed[1443],seed[658],seed[1630],seed[3514],seed[1902],seed[3293],seed[735],seed[358],seed[2478],seed[2712],seed[134],seed[2454],seed[594],seed[616],seed[823],seed[3453],seed[2721],seed[1076],seed[240],seed[3087],seed[245],seed[3943],seed[2370],seed[1842],seed[1394],seed[235],seed[1016],seed[2835],seed[1499],seed[839],seed[1371],seed[1083],seed[2713],seed[1217],seed[3213],seed[52],seed[3020],seed[2595],seed[292],seed[2710],seed[1921],seed[3341],seed[2338],seed[3487],seed[1939],seed[1418],seed[2983],seed[1723],seed[3634],seed[2599],seed[2376],seed[907],seed[3068],seed[2450],seed[1],seed[2992],seed[1693],seed[971],seed[2046],seed[3081],seed[1574],seed[1960],seed[572],seed[2510],seed[1234],seed[2700],seed[3246],seed[2501],seed[996],seed[1620],seed[3833],seed[795],seed[2685],seed[2277],seed[1513],seed[331],seed[2893],seed[3553],seed[1552],seed[1085],seed[3321],seed[3694],seed[3920],seed[480],seed[1179],seed[3198],seed[2896],seed[1141],seed[1634],seed[1763],seed[3295],seed[3623],seed[3248],seed[1216],seed[3057],seed[3245],seed[3366],seed[3123],seed[1661],seed[1260],seed[2041],seed[1088],seed[3599],seed[1629],seed[1377],seed[3436],seed[843],seed[2653],seed[813],seed[577],seed[283],seed[1832],seed[1953],seed[1241],seed[3191],seed[3380],seed[169],seed[3107],seed[2632],seed[320],seed[319],seed[1212],seed[2465],seed[448],seed[3834],seed[386],seed[355],seed[2076],seed[1649],seed[187],seed[3600],seed[615],seed[3700],seed[1163],seed[809],seed[2932],seed[1290],seed[863],seed[1884],seed[3573],seed[3438],seed[2590],seed[2437],seed[3825],seed[2611],seed[433],seed[645],seed[2011],seed[1906],seed[3182],seed[992],seed[2789],seed[598],seed[3095],seed[2631],seed[3252],seed[546],seed[2408],seed[3103],seed[2689],seed[2593],seed[2864],seed[623],seed[374],seed[3740],seed[2645],seed[1969],seed[3194],seed[1797],seed[1904],seed[3337],seed[3986],seed[3729],seed[47],seed[1640],seed[683],seed[3645],seed[1783],seed[3124],seed[1400],seed[3406],seed[197],seed[3203],seed[860],seed[833],seed[1295],seed[1536],seed[3186],seed[3806],seed[1828],seed[2616],seed[669],seed[2891],seed[3154],seed[3202],seed[470],seed[956],seed[89],seed[2899],seed[2609],seed[2324],seed[2826],seed[2387],seed[2898],seed[291],seed[941],seed[3746],seed[1456],seed[2317],seed[378],seed[2843],seed[444],seed[3327],seed[2206],seed[3995],seed[3728],seed[3403],seed[504],seed[3660],seed[620],seed[1314],seed[1778],seed[2777],seed[4015],seed[80],seed[2039],seed[1350],seed[3596],seed[724],seed[634],seed[2486],seed[41],seed[1081],seed[2459],seed[3965],seed[2068],seed[1857],seed[2005],seed[2065],seed[2259],seed[1809],seed[1202],seed[2538],seed[446],seed[1045],seed[429],seed[1249],seed[2544],seed[557],seed[2725],seed[902],seed[611],seed[1301],seed[2568],seed[2736],seed[1987],seed[832],seed[394],seed[1342],seed[3249],seed[2037],seed[1364],seed[2944],seed[2796],seed[224],seed[1027],seed[553],seed[2563],seed[1633],seed[3157],seed[3592],seed[1345],seed[2180],seed[1937],seed[2456],seed[2714],seed[2435],seed[2352],seed[3538],seed[533],seed[2771],seed[322],seed[2167],seed[1066],seed[438],seed[3882],seed[3537],seed[2995],seed[1541],seed[227],seed[2288],seed[3268],seed[827],seed[3666],seed[1005],seed[1341],seed[1127],seed[3723],seed[299],seed[753],seed[702],seed[2402],seed[1022],seed[1266],seed[481],seed[899],seed[3021],seed[2901],seed[1907],seed[259],seed[1340],seed[1180],seed[2060],seed[1830],seed[2168],seed[329],seed[1720],seed[68],seed[2702],seed[1185],seed[1835],seed[3361],seed[464],seed[3783],seed[3110],seed[3849],seed[3368],seed[37],seed[3513],seed[581],seed[749],seed[2149],seed[2910],seed[3846],seed[3784],seed[2102],seed[2426],seed[3927],seed[1467],seed[1475],seed[3437],seed[432],seed[401],seed[2764],seed[368],seed[309],seed[3836],seed[3713],seed[1654],seed[59],seed[97],seed[3083],seed[1892],seed[2745],seed[1518],seed[3650],seed[2131],seed[457],seed[2682],seed[3025],seed[3479],seed[1671],seed[2489],seed[77],seed[2112],seed[2344],seed[711],seed[2760],seed[1507],seed[1911],seed[3359],seed[3102],seed[2043],seed[3747],seed[391],seed[3942],seed[3072],seed[1426],seed[1235],seed[697],seed[1806],seed[2358],seed[3490],seed[915],seed[258],seed[1200],seed[2868],seed[1148],seed[1437],seed[1511],seed[514],seed[2455],seed[417],seed[877],seed[1041],seed[177],seed[2583],seed[788],seed[1227],seed[3674],seed[1665],seed[1867],seed[2844],seed[2951],seed[3775],seed[1190],seed[1698],seed[2965],seed[127],seed[1001],seed[3510],seed[3008],seed[3715],seed[2770],seed[4065],seed[145],seed[1936],seed[869],seed[151],seed[3903],seed[1749],seed[1846],seed[2798],seed[492],seed[2430],seed[844],seed[495],seed[800],seed[910],seed[3506],seed[1674],seed[2812],seed[3096],seed[969],seed[2743],seed[3050],seed[857],seed[1033],seed[663],seed[3693],seed[3063],seed[155],seed[2164],seed[1169],seed[1356],seed[3261],seed[1450],seed[3497],seed[2418],seed[2850],seed[50],seed[2117],seed[4039],seed[3758],seed[1877],seed[1715],seed[324],seed[972],seed[1645],seed[1178],seed[373],seed[1488],seed[3048],seed[2055],seed[1427],seed[26],seed[379],seed[808],seed[1440],seed[4084],seed[2421],seed[1140],seed[2976],seed[3823],seed[2559],seed[3522],seed[2640],seed[1868],seed[2818],seed[3016],seed[3176],seed[1900],seed[478],seed[654],seed[1370],seed[1714],seed[3821],seed[1412],seed[3980],seed[3452],seed[2988],seed[1113],seed[3710],seed[786],seed[649],seed[3333],seed[4080],seed[883],seed[2283],seed[1932],seed[3854],seed[1922],seed[3706],seed[3212],seed[3099],seed[1143],seed[3085],seed[629],seed[842],seed[3101],seed[3868],seed[1927],seed[961],seed[2364],seed[2495],seed[3983],seed[86],seed[3256],seed[2423],seed[3638],seed[4041],seed[1390],seed[252],seed[1871],seed[1259],seed[1847],seed[4030],seed[1648],seed[342],seed[2542],seed[655],seed[878],seed[2786],seed[3384],seed[3552],seed[3891],seed[1431],seed[2212],seed[1455],seed[1878],seed[300],seed[2639],seed[2614],seed[3350],seed[3168],seed[2116],seed[2572],seed[1554],seed[1108],seed[3483],seed[3221],seed[203],seed[1478],seed[92],seed[950],seed[1553],seed[3851],seed[1062],seed[387],seed[787],seed[1012],seed[1726],seed[2329],seed[3736],seed[1274],seed[3496],seed[3367],seed[726],seed[3717],seed[3754],seed[1053],seed[3652],seed[1616],seed[424],seed[3211],seed[419],seed[2792],seed[1524],seed[3024],seed[503],seed[3431],seed[276],seed[1192],seed[2851],seed[2819],seed[2558],seed[3542],seed[3533],seed[3201],seed[137],seed[2494],seed[1373],seed[2741],seed[36],seed[3056],seed[2986],seed[2309],seed[399],seed[390],seed[867],seed[3764],seed[2555],seed[3108],seed[213],seed[2357],seed[2445],seed[2902],seed[2781],seed[2363],seed[3074],seed[2340],seed[761],seed[2513],seed[2040],seed[1718],seed[3789],seed[229],seed[1395],seed[2929],seed[2575],seed[3343],seed[2954],seed[1941],seed[855],seed[3826],seed[3940],seed[678],seed[2442],seed[3465],seed[3036],seed[3689],seed[2610],seed[696],seed[3730],seed[3287],seed[436],seed[2017],seed[2030],seed[549],seed[816],seed[2657],seed[3861],seed[1568],seed[1562],seed[434],seed[2135],seed[1592],seed[2401],seed[251],seed[2356],seed[1705],seed[376],seed[306],seed[2215],seed[2726],seed[2477],seed[3028],seed[3714],seed[1287],seed[1311],seed[3267],seed[274],seed[1430],seed[226],seed[2010],seed[502],seed[1482],seed[991],seed[2160],seed[610],seed[3504],seed[2293],seed[3997],seed[260],seed[1759],seed[3755],seed[3489],seed[1560],seed[3263],seed[173],seed[2140],seed[1285],seed[2587],seed[801],seed[2471],seed[1545],seed[2950],seed[273],seed[635],seed[35],seed[3111],seed[363],seed[2388],seed[3531],seed[3773],seed[2110],seed[241],seed[3117],seed[1897],seed[2779],seed[427],seed[3400],seed[687],seed[1767],seed[1193],seed[569],seed[2382],seed[2330],seed[794],seed[3372],seed[785],seed[1746],seed[681],seed[3984],seed[3896],seed[3901],seed[3994],seed[1567],seed[1044],seed[3079],seed[325],seed[2534],seed[1619],seed[1711],seed[1879],seed[326],seed[2553],seed[1232],seed[1751],seed[2748],seed[952],seed[483],seed[819],seed[507],seed[2057],seed[79],seed[2020],seed[1451],seed[1777],seed[2093],seed[1245],seed[1849],seed[776],seed[3898],seed[2084],seed[3273],seed[876],seed[738],seed[1191],seed[354],seed[1901],seed[2451],seed[804],seed[3325],seed[1396],seed[76],seed[3549],seed[3187],seed[2487],seed[1840],seed[3047],seed[2620],seed[1942],seed[4078],seed[3532],seed[1547],seed[4024],seed[614],seed[922],seed[2801],seed[3105],seed[2564],seed[2841],seed[3338],seed[3760],seed[2424],seed[817],seed[1258],seed[1078],seed[3466],seed[3576],seed[1461],seed[1300],seed[186],seed[1925],seed[3907],seed[3462],seed[163],seed[2808],seed[330],seed[798],seed[3291],seed[803],seed[3708],seed[3336],seed[2696],seed[1402],seed[3525],seed[3979],seed[3671],seed[3850],seed[183],seed[1933],seed[1952],seed[2541],seed[2342],seed[2622],seed[2594],seed[3259],seed[695],seed[1335],seed[2213],seed[2145],seed[2848],seed[1521],seed[3864],seed[3423],seed[1292],seed[2322],seed[1152],seed[2753],seed[1470],seed[987],seed[3751],seed[411],seed[1065],seed[345],seed[1793],seed[1291],seed[1293],seed[2222],seed[2884],seed[2975],seed[2443],seed[3383],seed[2768],seed[2049],seed[3053],seed[1247],seed[1404],seed[3551],seed[590],seed[831],seed[506],seed[409],seed[1406],seed[3495],seed[3686],seed[555],seed[1358],seed[4082],seed[1220],seed[1151],seed[344],seed[2158],seed[78],seed[1142],seed[4068],seed[2514],seed[2263],seed[754],seed[375],seed[3209],seed[1063],seed[1176],seed[1584],seed[1423],seed[449],seed[3315],seed[208],seed[2059],seed[3842],seed[1347],seed[3316],seed[3439],seed[2069],seed[2822],seed[3470],seed[102],seed[249],seed[541],seed[3426],seed[3961],seed[1319],seed[3445],seed[2304],seed[1570],seed[3344],seed[3559],seed[2272],seed[2407],seed[1360],seed[1004],seed[2678],seed[262],seed[1731],seed[3948],seed[1614],seed[2927],seed[3142],seed[1020],seed[2464],seed[1339],seed[2968],seed[3857],seed[1174],seed[4056],seed[4036],seed[2268],seed[136],seed[1155],seed[3370],seed[742],seed[2674],seed[3322],seed[743],seed[712],seed[4061],seed[2809],seed[1559],seed[1557],seed[3217],seed[2044],seed[3032],seed[1336],seed[362],seed[3697],seed[1975],seed[1949],seed[2229],seed[2378],seed[2075],seed[980],seed[3779],seed[3014],seed[2007],seed[3695],seed[3603],seed[3923],seed[2663],seed[1317],seed[3459],seed[1946],seed[3547],seed[3109],seed[195],seed[3238],seed[2284],seed[1401],seed[2498],seed[1851],seed[3262],seed[2091],seed[2087],seed[3681],seed[731],seed[10],seed[201],seed[1608],seed[1866],seed[2739],seed[2990],seed[2279],seed[2249],seed[3739],seed[2207],seed[1821],seed[3141],seed[2500],seed[3241],seed[4025],seed[2719],seed[315],seed[3702],seed[1031],seed[3448],seed[1189],seed[3369],seed[3159],seed[3144],seed[3976],seed[3959],seed[3737],seed[1954],seed[1253],seed[3118],seed[3752],seed[2452],seed[1156],seed[1701],seed[2473],seed[191],seed[2174],seed[3772],seed[3523],seed[165],seed[3],seed[2188],seed[1374],seed[2876],seed[3974],seed[3519],seed[3945],seed[2603],seed[2939],seed[3545],seed[912],seed[565],seed[184],seed[1566],seed[1091],seed[2890],seed[1918],seed[1346],seed[1745],seed[3482],seed[2348],seed[3933],seed[3738],seed[2275],seed[1898],seed[2225],seed[667],seed[3092],seed[2612],seed[3193],seed[672],seed[474],seed[1117],seed[830],seed[3023],seed[3967],seed[2061],seed[3416],seed[494],seed[54],seed[3711],seed[3804],seed[1772],seed[1188],seed[2925],seed[2208],seed[1721],seed[3051],seed[3152],seed[3800],seed[2144],seed[1860],seed[2391],seed[3289],seed[1165],seed[3631],seed[289],seed[3769],seed[232],seed[3848],seed[2775],seed[2856],seed[3210],seed[2281],seed[2729],seed[1989],seed[686],seed[605],seed[600],seed[296],seed[706],seed[1514],seed[1029],seed[2744],seed[2148],seed[1221],seed[2336],seed[3376],seed[48],seed[435],seed[179],seed[2232],seed[450],seed[222],seed[2546],seed[3323],seed[3451],seed[1785],seed[895],seed[2987],seed[3420],seed[3763],seed[1248],seed[3546],seed[3319],seed[234],seed[2171],seed[2032],seed[2852],seed[1818],seed[3892],seed[3735],seed[2815],seed[2214],seed[3869],seed[880],seed[293],seed[4049],seed[908],seed[3388],seed[23],seed[193],seed[3398],seed[2367],seed[2785],seed[2062],seed[2832],seed[2875],seed[684],seed[1534],seed[2374],seed[2977],seed[1298],seed[3741],seed[3993],seed[990],seed[2080],seed[2972],seed[3039],seed[1869],seed[3937],seed[722],seed[3133],seed[2313],seed[1862],seed[2924],seed[556],seed[3455],seed[1573],seed[1479],seed[1637],seed[1760],seed[3175],seed[2961],seed[2012],seed[1223],seed[56],seed[2897],seed[2958],seed[141],seed[641],seed[2776],seed[679],seed[3204],seed[2916],seed[1623],seed[624],seed[6],seed[1606],seed[887],seed[2441],seed[2203],seed[491],seed[31],seed[3687],seed[886],seed[118],seed[2695],seed[1369],seed[242],seed[341],seed[2429],seed[736],seed[81],seed[217],seed[2349],seed[285],seed[3947],seed[3064],seed[847],seed[2940],seed[1702],seed[1983],seed[4053],seed[1409],seed[2077],seed[3831],seed[2125],seed[57],seed[2694],seed[1825],seed[1587],seed[3958],seed[905],seed[1469],seed[1145],seed[1146],seed[3254],seed[58],seed[2254],seed[1484],seed[935],seed[625],seed[3872],seed[3243],seed[3704],seed[2150],seed[659],seed[2787],seed[1366],seed[3679],seed[796],seed[1262],seed[3795],seed[1526],seed[3391],seed[2209],seed[2720],seed[1415],seed[3399],seed[2183],seed[909],seed[3893],seed[2094],seed[3557],seed[115],seed[3169],seed[3362],seed[3575],seed[1361],seed[160],seed[3279],seed[2874],seed[1986],seed[1264],seed[2579],seed[4066],seed[542],seed[3748],seed[2172],seed[1037],seed[1889],seed[496],seed[2921],seed[1457],seed[3707],seed[3585],seed[124],seed[2205],seed[778],seed[1905],seed[874],seed[1811],seed[1981],seed[3765],seed[2413],seed[2946],seed[3996],seed[3624],seed[3879],seed[4020],seed[1182],seed[1125],seed[1422],seed[1057],seed[1104],seed[1399],seed[3146],seed[951],seed[236],seed[476],seed[1102],seed[428],seed[3598],seed[1742],seed[2806],seed[2831],seed[1870],seed[2053],seed[2347],seed[871],seed[2202],seed[793],seed[1489],seed[4021],seed[3234],seed[1713],seed[488],seed[3125],seed[3955],seed[3314],seed[2731],seed[2833],seed[2325],seed[3132],seed[2918],seed[2056],seed[287],seed[1666],seed[2492],seed[396],seed[1873],seed[1320],seed[1709],seed[2701],seed[2982],seed[1957],seed[51],seed[824],seed[2434],seed[1080],seed[2189],seed[270],seed[2107],seed[21],seed[692],seed[67],seed[3460],seed[3017],seed[1744],seed[2545],seed[1845],seed[810],seed[1011],seed[2754],seed[527],seed[228],seed[1914],seed[2051],seed[3544],seed[2854],seed[3253],seed[1122],seed[834],seed[462],seed[152],seed[1795],seed[3956],seed[1173],seed[1284],seed[465],seed[1669],seed[1678],seed[3724],seed[3574],seed[3633],seed[812],seed[340],seed[1222],seed[946],seed[2462],seed[3389],seed[2591],seed[660],seed[3621],seed[2634],seed[243],seed[3616],seed[1736],seed[562],seed[1046],seed[3508],seed[2190],seed[117],seed[3662],seed[1071],seed[1302],seed[3517],seed[2532],seed[2409],seed[2200],seed[214],seed[1392],seed[3651],seed[1815],seed[3000],seed[1114],seed[2292],seed[1881],seed[2438],seed[1627],seed[1271],seed[3790],seed[1943],seed[2031],seed[1106],seed[1454],seed[2613],seed[3290],seed[894],seed[1908],seed[3299],seed[101],seed[2238],seed[3541],seed[1228],seed[646],seed[2960],seed[1299],seed[936],seed[32],seed[3353],seed[3818],seed[369],seed[2879],seed[1225],seed[2684],seed[756],seed[1378],seed[311],seed[2377],seed[2375],seed[3529],seed[1580],seed[2446],seed[1564],seed[3918],seed[2196],seed[2396],seed[458],seed[1150],seed[1948],seed[64],seed[1230],seed[962],seed[937],seed[3719],seed[18],seed[2319],seed[2919],seed[2416],seed[602],seed[917],seed[3145],seed[1441],seed[3358],seed[2767],seed[2993],seed[3954],seed[2386],seed[2226],seed[3410],seed[3811],seed[2499],seed[1915],seed[400],seed[3292],seed[3564],seed[3224],seed[1313],seed[3649],seed[2153],seed[1931],seed[913],seed[3718],seed[3059],seed[747],seed[975],seed[2882],seed[3759],seed[1602],seed[3022],seed[1556],seed[901],seed[1509],seed[2649],seed[2311],seed[1432],seed[1330],seed[1730],seed[680],seed[3692],seed[560],seed[3480],seed[3664],seed[1756],seed[2070],seed[2333],seed[3609],seed[3659],seed[212],seed[1413],seed[573],seed[2233],seed[1307],seed[1375],seed[2035],seed[3356],seed[2855],seed[156],seed[1681],seed[1238],seed[4042],seed[1231],seed[3632],seed[2381],seed[2550],seed[2635],seed[3771],seed[3732],seed[467],seed[159],seed[3340],seed[3870],seed[2242],seed[1382],seed[2949],seed[3060],seed[132],seed[441],seed[1644],seed[1612],seed[2025],seed[1407],seed[642],seed[2569],seed[3647],seed[4064],seed[11],seed[2504],seed[1069],seed[1486],seed[3414],seed[2525],seed[2166],seed[1344],seed[2920],seed[2425],seed[3843],seed[1476],seed[3121],seed[1015],seed[1119],seed[3113],seed[2655],seed[38],seed[2024],seed[2294],seed[3478],seed[412],seed[1647],seed[1211],seed[70],seed[526],seed[2942],seed[1471],seed[1343],seed[1993],seed[3345],seed[3819],seed[1097],seed[1021],seed[3932],seed[2727],seed[456],seed[1517],seed[3677],seed[3467],seed[13],seed[1532],seed[700],seed[3646],seed[3239],seed[269],seed[1105],seed[317],seed[561],seed[1690],seed[1028],seed[3231],seed[558],seed[3371],seed[3163],seed[1408],seed[1003],seed[2469],seed[205],seed[3881],seed[1646],seed[4008],seed[1017],seed[2804],seed[2524],seed[1226],seed[1968],seed[2643],seed[1675],seed[202],seed[3427],seed[1095],seed[1662],seed[2857],seed[1595],seed[24],seed[1160],seed[85],seed[885],seed[1495],seed[2605],seed[1970],seed[882],seed[2650],seed[791],seed[3257],seed[2570],seed[889],seed[925],seed[2888],seed[3306],seed[3071],seed[2173],seed[3844],seed[3463],seed[1158],seed[3309],seed[1657],seed[2554],seed[295],seed[1326],seed[2157],seed[334],seed[2165],seed[3046],seed[892],seed[3173],seed[1333],seed[499],seed[1880],seed[3419],seed[279],seed[3461],seed[918],seed[72],seed[3320],seed[3781],seed[931],seed[2991],seed[1635],seed[3225],seed[2320],seed[2585],seed[1782],seed[377],seed[3762],seed[4011],seed[775],seed[3630],seed[4083],seed[2562],seed[1239],seed[3223],seed[2926],seed[701],seed[1244],seed[1072],seed[1208],seed[1490],seed[290],seed[1137],seed[4028],seed[989],seed[1459],seed[3318],seed[1773],seed[53],seed[636],seed[1572],seed[1492],seed[1420],seed[3563],seed[3999],seed[2006],seed[1590],seed[2406],seed[4022],seed[1010],seed[1162],seed[1836],seed[3015],seed[675],seed[3805],seed[508],seed[2820],seed[3502],seed[2783],seed[3250],seed[1498],seed[49],seed[1824],seed[2088],seed[1254],seed[1079],seed[2565],seed[43],seed[699],seed[3526],seed[2072],seed[845],seed[3283],seed[2703],seed[1306],seed[1727],seed[3527],seed[2512],seed[1099],seed[1483],seed[2606],seed[1294],seed[767],seed[4050],seed[1965],seed[997],seed[1296],seed[1448],seed[1466],seed[1205],seed[1309],seed[613],seed[668],seed[1875],seed[691],seed[4069],seed[2089],seed[3591],seed[3981],seed[3982],seed[530],seed[73],seed[1485],seed[3192],seed[1844],seed[162],seed[3165],seed[1329],seed[1741],seed[3683],seed[576],seed[2625],seed[3776],seed[17],seed[3709],seed[1684],seed[1438],seed[1136],seed[1365],seed[1955],seed[622],seed[1118],seed[1243],seed[402],seed[1058],seed[2228],seed[3242],seed[1978],seed[178],seed[2668],seed[3200],seed[911],seed[3890],seed[2706],seed[3571],seed[1397],seed[2536],seed[3150],seed[2461],seed[482],seed[2104],seed[534],seed[2581],seed[4072],seed[2318],seed[2314],seed[1529],seed[3301],seed[1039],seed[868],seed[3127],seed[3528],seed[1376],seed[1679],seed[3422],seed[3579],seed[4038],seed[2989],seed[3106],seed[579],seed[3317],seed[3636],seed[1052],seed[3911],seed[257],seed[1909],seed[853],seed[2661],seed[2795],seed[3876],seed[2432],seed[2139],seed[1446],seed[677],seed[2734],seed[2828],seed[4044],seed[3001],seed[1372],seed[2118],seed[765],seed[254],seed[3619],seed[2930],seed[1683],seed[3815],seed[1694],seed[3382],seed[963],seed[2911],seed[4043],seed[19],seed[2170],seed[1428],seed[1515],seed[3595],seed[861],seed[280],seed[1996],seed[3364],seed[3185],seed[2521],seed[3886],seed[2194],seed[3499],seed[2970],seed[741],seed[2704],seed[571],seed[218],seed[1754],seed[1753],seed[1589],seed[3147],seed[2759],seed[3897],seed[3005],seed[2578],seed[1770],seed[2267],seed[2101],seed[954],seed[2355],seed[2129],seed[1281],seed[2155],seed[688],seed[28],seed[4074],seed[1823],seed[2136],seed[671],seed[1398],seed[1391],seed[1883],seed[2629],seed[717],seed[1591],seed[1184],seed[897],seed[140],seed[1839],seed[627],seed[3614],seed[2866],seed[1135],seed[2867],seed[3026],seed[1194],seed[442],seed[1807],seed[750],seed[3569],seed[1579],seed[1771],seed[1077],seed[2733],seed[238],seed[2475],seed[626],seed[2909],seed[693],seed[2193],seed[2842],seed[3172],seed[3511],seed[548],seed[4060],seed[1703],seed[3442],seed[2711],seed[3908],seed[1009],seed[3164],seed[2191],seed[2531],seed[256],seed[4077],seed[3031],seed[2305],seed[3076],seed[705],seed[942],seed[3884],seed[119],seed[1963],seed[3251],seed[2551],seed[196],seed[2241],seed[3644],seed[1596],seed[888],seed[1363],seed[2906],seed[168],seed[61],seed[944],seed[2738],seed[815],seed[353],seed[490],seed[420],seed[2933],seed[107],seed[1442],seed[3678],seed[3394],seed[209],seed[593],seed[2928],seed[188],seed[1318],seed[3395],seed[3417],seed[2935],seed[2015],seed[3970],seed[998],seed[837],seed[263],seed[799],seed[2580],seed[2162],seed[3612],seed[2732],seed[498],seed[2085],seed[2253],seed[339],seed[1387],seed[2889],seed[1765],seed[1133],seed[2098],seed[2752],seed[923],seed[2127],seed[3313],seed[3434],seed[367],seed[924],seed[323],seed[2788],seed[3122],seed[485],seed[2197],seed[3568],seed[2398],seed[1973],seed[2114],seed[380],seed[3007],seed[2286],seed[3070],seed[1103],seed[740],seed[2519],seed[3975],seed[575],seed[719],seed[2236],seed[780],seed[1600],seed[3924],seed[2100],seed[3255],seed[2250],seed[2664],seed[2937],seed[1604],seed[1935],seed[708],seed[3062],seed[2244],seed[566],seed[1837],seed[1240],seed[1977],seed[1601],seed[1940],seed[3653],seed[698],seed[154],seed[3658],seed[3216],seed[505],seed[729],seed[1452],seed[3035],seed[1658],seed[2862],seed[1123],seed[2681],seed[3774],seed[3274],seed[1171],seed[3003],seed[9],seed[3390],seed[835],seed[981],seed[2686],seed[2677],seed[2608],seed[1138],seed[884],seed[2567],seed[2496],seed[4091],seed[1872],seed[2886],seed[3605],seed[1279],seed[2626],seed[966],seed[3867],seed[3112],seed[3349],seed[2028],seed[2397],seed[2747],seed[587],seed[430],seed[2474],seed[1084],seed[3909],seed[2237],seed[519],seed[3566],seed[2296],seed[100],seed[2383],seed[3377],seed[303],seed[3027],seed[1789],seed[1530],seed[1368],seed[3668],seed[3138],seed[2953],seed[3757],seed[25],seed[2662],seed[3272],seed[1512],seed[305],seed[3428],seed[3550],seed[3657],seed[1491],seed[4058],seed[327],seed[3180],seed[3304],seed[2830],seed[858],seed[960],seed[2627],seed[3565],seed[2248],seed[189],seed[2334],seed[2637],seed[2604],seed[2883],seed[3828],seed[4023],seed[2887],seed[133],seed[343],seed[3931],seed[2354],seed[1013],seed[2530],seed[3114],seed[2628],seed[4095],seed[580],seed[2332],seed[3900],seed[3196],seed[1668],seed[1000],seed[93],seed[1653],seed[1269],seed[45],seed[720],seed[1094],seed[2130],seed[3935],seed[2054],seed[1859],seed[393],seed[1324],seed[1740],seed[3207],seed[1739],seed[4094],seed[2493],seed[3094],seed[2769],seed[2692],seed[1689],seed[298],seed[233],seed[3562],seed[1819],seed[250],seed[2722],seed[103],seed[170],seed[2186],seed[2617],seed[3044],seed[1075],seed[515],seed[985],seed[2063],seed[2638],seed[2086],seed[2274],seed[940],seed[520],seed[4040],seed[3602],seed[1332],seed[1700],seed[2724],seed[2224],seed[1788],seed[1101],seed[3570],seed[2204],seed[2966],seed[3780],seed[3750],seed[3435],seed[545],seed[1331],seed[1256],seed[1038],seed[1947],seed[1073],seed[3174],seed[2278],seed[2756],seed[1733],seed[3663],seed[1886],seed[2428],seed[1074],seed[1801],seed[3220],seed[2824],seed[484],seed[2103],seed[4027],seed[3019],seed[3458],seed[852],seed[1747],seed[2900],seed[2520],seed[866],seed[967],seed[570],seed[1445],seed[900],seed[2528],seed[1502],seed[2690],seed[1018],seed[1803],seed[207],seed[1110],seed[1494],seed[4018],seed[1187],seed[930],seed[811],seed[3934],seed[3135],seed[948],seed[955],seed[1656],seed[3930],seed[142],seed[1799],seed[1798],seed[1991],seed[609],seed[725],seed[2351],seed[451],seed[46],seed[893],seed[2589],seed[3796],seed[1791],seed[3066],seed[1691],seed[3838],seed[3247],seed[1334],seed[974],seed[1643],seed[596],seed[2109],seed[510],seed[559],seed[3342],seed[2652],seed[2050],seed[225],seed[4033],seed[1548],seed[1535],seed[445],seed[3346],seed[1435],seed[1276],seed[820],seed[2300],seed[3149],seed[3847],seed[3643],seed[2517],seed[982],seed[2303],seed[1167],seed[657],seed[3987],seed[1393],seed[1642],seed[2871],seed[4063],seed[2647],seed[1899],seed[2509],seed[199],seed[3871],seed[3964],seed[172],seed[770],seed[739],seed[497],seed[3797],seed[1813],seed[2790],seed[1047],seed[3407],seed[3311],seed[523],seed[1651],seed[3807],seed[589],seed[2584],seed[3661],seed[1624],seed[1323],seed[3885],seed[2751],seed[1796],seed[2914],seed[1060],seed[200],seed[976],seed[3120],seed[2680],seed[732],seed[3977],seed[2247],seed[1107],seed[2648],seed[2936],seed[1050],seed[1923],seed[2192],seed[1603],seed[74],seed[42],seed[486],seed[3782],seed[1019],seed[1421],seed[1885],seed[2199],seed[2586],seed[3137],seed[3904],seed[1115],seed[1149],seed[106],seed[3441],seed[2540],seed[3468],seed[2847],seed[1810],seed[2415],seed[2705],seed[318],seed[2571],seed[2122],seed[346],seed[2400],seed[3720],seed[3214],seed[2757],seed[2894],seed[3827],seed[1381],seed[2152],seed[2252],seed[3115],seed[2548],seed[734],seed[1976],seed[372],seed[16],seed[3922],seed[3655],seed[2723],seed[466],seed[947],seed[619],seed[3091],seed[2384],seed[1834],seed[335],seed[1132],seed[422],seed[1035],seed[447],seed[2380],seed[1168],seed[792],seed[2597],seed[4087],seed[153],seed[516],seed[3509],seed[3852],seed[113],seed[3156],seed[2908],seed[715],seed[87],seed[2913],seed[2881],seed[1628],seed[469],seed[1116],seed[1519],seed[1650],seed[314],seed[1425],seed[1386],seed[2353],seed[763],seed[3012],seed[1664],seed[2147],seed[3963],seed[3587],seed[1577],seed[2800],seed[755],seed[2687],seed[2310],seed[3088],seed[3808],seed[1082],seed[512],seed[4093],seed[1261],seed[1750],seed[1586],seed[584],seed[164],seed[3770],seed[3586],seed[2817],seed[3421],seed[1453],seed[2346],seed[585],seed[2485],seed[760],seed[403],seed[359],seed[1447],seed[2036],seed[2276],seed[3183],seed[2002],seed[2295],seed[4086],seed[1025],seed[2120],seed[551],seed[779],seed[1542],seed[3043],seed[3171],seed[3303],seed[2598],seed[3731],seed[2577],seed[2411],seed[3915],seed[1990],seed[3648],seed[2892],seed[1338],seed[1242],seed[3244],seed[3049],seed[2903],seed[3086],seed[2337],seed[1626],seed[906],seed[2182],seed[653],seed[3433],seed[371],seed[821],seed[55],seed[2742],seed[1195],seed[1636],seed[3676],seed[2113],seed[864],seed[3312],seed[3803],seed[1144],seed[3613],seed[398],seed[4029],seed[2071],seed[4055],seed[210],seed[2027],seed[1516],seed[2359],seed[1578],seed[1051],seed[261],seed[1219],seed[3424],seed[3179],seed[1800],seed[3953],seed[2688],seed[3874],seed[3494],seed[3601],seed[3412],seed[22],seed[768],seed[1549],seed[2312],seed[1894],seed[1067],seed[1555],seed[3045],seed[1615],seed[1599],seed[1109],seed[673],seed[1569],seed[3902],seed[88],seed[532],seed[146],seed[366],seed[221],seed[479],seed[3310],seed[3578],seed[3227],seed[2003],seed[2985],seed[4054],seed[2014],seed[392],seed[814],seed[2670],seed[547],seed[487],seed[489],seed[977],seed[2774],seed[1233],seed[2772],seed[3802],seed[333],seed[1086],seed[360],seed[1098],seed[3308],seed[3073],seed[3627],seed[144],seed[2126],seed[986],seed[2019],seed[1699],seed[2405],seed[1315],seed[408],seed[1697],seed[1980],seed[2097],seed[348],seed[3703],seed[1768],seed[968],seed[3334],seed[3939],seed[3042],seed[2766],seed[3139],seed[2557],seed[1728],seed[2917],seed[1865],seed[3503],seed[3793],seed[2675],seed[1463],seed[1157],seed[1575],seed[2273],seed[1757],seed[1056],seed[255],seed[3286],seed[71],seed[123],seed[2730],seed[929],seed[1449],seed[3277],seed[524],seed[2285],seed[3957],seed[108],seed[3588],seed[1582],seed[150],seed[4046],seed[1288],seed[3457],seed[3691],seed[3926],seed[2878],seed[3866],seed[2301],seed[3929],seed[95],seed[1958],seed[30],seed[223],seed[599],seed[3787],seed[752],seed[2676],seed[2860],seed[3938],seed[3534],seed[2201],seed[62],seed[2042],seed[3298],seed[1561],seed[1474],seed[3829],seed[3197],seed[2588],seed[3498],seed[310],seed[781],seed[2410],seed[3799],seed[1995],seed[3583],seed[39],seed[2389],seed[710],seed[3788],seed[2912],seed[2811],seed[2266],seed[841],seed[2184],seed[2137],seed[2251],seed[397],seed[2083],seed[415],seed[3447],seed[3129],seed[3742],seed[220],seed[3604],seed[216],seed[468],seed[2161],seed[3734],seed[3222],seed[2502],seed[1214],seed[1852],seed[3500],seed[2794],seed[66],seed[1362],seed[3543],seed[1808],seed[643],seed[3756],seed[3328],seed[618],seed[2483],seed[2264],seed[2573],seed[662],seed[1804],seed[2394],seed[1916],seed[3034],seed[1403],seed[338],seed[875],seed[1738],seed[849],seed[1831],seed[3906],seed[3002],seed[586],seed[2582],seed[3488],seed[2243],seed[933],seed[3375],seed[1460],seed[63],seed[1717],seed[854],seed[2671],seed[957],seed[15],seed[3985],seed[773],seed[1439],seed[1994],seed[1988],seed[1890],seed[2282],seed[1111],seed[2073],seed[1410],seed[3794],seed[3952],seed[1436],seed[1054],seed[1966],seed[4034],seed[2735],seed[1351],seed[1673],seed[3998],seed[1480],seed[1280],seed[2636],seed[2302],seed[3916],seed[766],seed[3232],seed[3331],seed[1093],seed[1325],seed[2009],seed[2945],seed[198],seed[370],seed[1934],seed[443],seed[1609],seed[1354],seed[3469],seed[304],seed[336],seed[138],seed[1639],seed[789],seed[416],seed[3491],seed[2641],seed[943],seed[1388],seed[2576],seed[2984],seed[3348],seed[3443],seed[4071],seed[2082],seed[1695],seed[3656],seed[1638],seed[1252],seed[3128],seed[3669],seed[3476],seed[988],seed[2045],seed[1096],seed[631],seed[685],seed[3512],seed[1583],seed[3233],seed[1385],seed[3950],seed[1417],seed[452],seed[128],seed[3010],seed[1175],seed[1780],seed[1776],seed[1164],seed[3905],seed[4079],seed[1864],seed[347],seed[3778],seed[139],seed[682],seed[2457],seed[807],seed[2805],seed[2299],seed[2840],seed[1196],seed[351],seed[1812],seed[2460],seed[111],seed[230],seed[1161],seed[694],seed[2998],seed[2642],seed[3265],seed[116],seed[3567],seed[1998],seed[630],seed[1667],seed[3151],seed[727],seed[301],seed[730],seed[3365],seed[3450],seed[2658],seed[1468],seed[3798],seed[3270],seed[1945],seed[1186],seed[1321],seed[1312],seed[2529],seed[2458],seed[1533],seed[194],seed[3363],seed[829],seed[475],seed[3518],seed[248],seed[405],seed[1204],seed[3625],seed[1210],seed[2240],seed[3177],seed[850],seed[2141],seed[4085],seed[3404],seed[3628],seed[2709],seed[2699],seed[1224],seed[578],seed[3743],seed[3877],seed[1631],seed[564],seed[535],seed[3440],seed[1967],seed[3925],seed[2621],seed[2797],seed[1962],seed[3167],seed[3078],seed[2959],seed[2829],seed[461],seed[3584],seed[2],seed[1303],seed[1500],seed[2623],seed[1607],seed[772],seed[862],seed[2837],seed[3786],seed[1893],seed[2096],seed[928],seed[3611],seed[1622],seed[1250],seed[1551],seed[3104],seed[1982],seed[525],seed[3093],seed[3622],seed[2799],seed[3392],seed[1613],seed[4062],seed[2934],seed[2869],seed[4076],seed[3184],seed[1197],seed[973],seed[3607],seed[246],seed[2466],seed[2872],seed[418],seed[3944],seed[2849],seed[2969],seed[2047],seed[2602],seed[2307],seed[356],seed[1748],seed[1672],seed[1049],seed[3582],seed[2343],seed[3004],seed[3520],seed[4081],seed[3858],seed[1755],seed[1289],seed[978],seed[1121],seed[970],seed[1429],seed[3084],seed[83],seed[1888],seed[1068],seed[2439],seed[2198],seed[337],seed[4089],seed[2269],seed[2372],seed[3266],seed[211],seed[190],seed[3968],seed[714],seed[1680],seed[4092],seed[282],seed[1030],seed[995],seed[539],seed[1652],seed[44],seed[2784],seed[2737],seed[3456],seed[999],seed[2646],seed[1297],seed[536],seed[3332],seed[1353],seed[1632],seed[192],seed[1272],seed[40],seed[3475],seed[2328],seed[4012],seed[1540],seed[2159],seed[2825],seed[3302],seed[4],seed[984],seed[1465],seed[1531],seed[3561],seed[3810],seed[1092],seed[3978],seed[582],seed[1971],seed[2185],seed[477],seed[1112],seed[4045],seed[472],seed[239],seed[473],seed[3832],seed[1383],seed[3733],seed[1305],seed[3134],seed[1896],seed[2339],seed[2067],seed[4004],seed[1024],seed[3912],seed[388],seed[2210],seed[2491],seed[3744],seed[3992],seed[2853],seed[2142],seed[1732],seed[3620],seed[316],seed[2099],seed[3887],seed[1206],seed[2938],seed[746],seed[2683],seed[3271],seed[1707],seed[2000],seed[891],seed[3880],seed[983],seed[650],seed[607],seed[3485],seed[2468],seed[1959],seed[2974],seed[2106],seed[674],seed[2216],seed[1929],seed[938],seed[4001],seed[3402],seed[3888],seed[2124],seed[2904],seed[4059],seed[2566],seed[994],seed[737],seed[3859],seed[3555],seed[3235],seed[608],seed[1611],seed[2119],seed[1621],seed[595],seed[2480],seed[540],seed[2260],seed[3722],seed[1563],seed[563],seed[2081],seed[1126],seed[4088],seed[1659],seed[1268],seed[2345],seed[1283],seed[1719],seed[3357],seed[644],seed[2708],seed[2802],seed[1685],seed[550],seed[1861],seed[2561],seed[3329],seed[3188],seed[1641],seed[2518],seed[439],seed[2026],seed[2331],seed[3535],seed[1040],seed[3530],seed[3385],seed[1558]}; 
//        seed15 <= {seed[603],seed[123],seed[592],seed[851],seed[4074],seed[928],seed[1023],seed[1200],seed[284],seed[1763],seed[566],seed[267],seed[1970],seed[3437],seed[3311],seed[1924],seed[476],seed[3329],seed[2712],seed[2040],seed[526],seed[3334],seed[1001],seed[3335],seed[1408],seed[1523],seed[1945],seed[4093],seed[2339],seed[1895],seed[536],seed[326],seed[887],seed[3034],seed[3885],seed[1885],seed[2805],seed[1343],seed[1144],seed[301],seed[2110],seed[2594],seed[3516],seed[354],seed[1624],seed[3195],seed[1540],seed[72],seed[2421],seed[1340],seed[3116],seed[1549],seed[2385],seed[1626],seed[425],seed[190],seed[1423],seed[2199],seed[1859],seed[1269],seed[1896],seed[1515],seed[2020],seed[3806],seed[4062],seed[1602],seed[1359],seed[938],seed[2679],seed[1092],seed[203],seed[909],seed[1564],seed[2830],seed[482],seed[1159],seed[561],seed[4083],seed[582],seed[2113],seed[389],seed[3048],seed[68],seed[3089],seed[2903],seed[2349],seed[74],seed[2999],seed[3562],seed[3032],seed[3825],seed[1630],seed[2327],seed[744],seed[3850],seed[2375],seed[819],seed[2478],seed[1411],seed[544],seed[4015],seed[2450],seed[3463],seed[1766],seed[2201],seed[455],seed[3384],seed[2939],seed[132],seed[3002],seed[438],seed[1548],seed[4005],seed[1258],seed[3213],seed[2891],seed[699],seed[1636],seed[332],seed[3628],seed[2657],seed[2489],seed[208],seed[325],seed[3888],seed[722],seed[2852],seed[2513],seed[2274],seed[1939],seed[3655],seed[1714],seed[2568],seed[2212],seed[2445],seed[1043],seed[3613],seed[569],seed[2119],seed[4077],seed[1476],seed[554],seed[3193],seed[3889],seed[3391],seed[1202],seed[4043],seed[2610],seed[3462],seed[4054],seed[2018],seed[1058],seed[1036],seed[2543],seed[3596],seed[1000],seed[992],seed[3529],seed[1363],seed[2909],seed[3151],seed[63],seed[3778],seed[3059],seed[3044],seed[1305],seed[1450],seed[3589],seed[1937],seed[172],seed[159],seed[487],seed[1510],seed[899],seed[3107],seed[3421],seed[1122],seed[491],seed[266],seed[2976],seed[146],seed[1274],seed[115],seed[1035],seed[2726],seed[1779],seed[1090],seed[3394],seed[3839],seed[1216],seed[783],seed[2943],seed[3216],seed[3840],seed[2207],seed[486],seed[3123],seed[1625],seed[1740],seed[2680],seed[3261],seed[937],seed[211],seed[2924],seed[794],seed[3077],seed[884],seed[4031],seed[3231],seed[2573],seed[2149],seed[3785],seed[117],seed[1662],seed[3570],seed[3648],seed[2325],seed[3924],seed[4010],seed[1977],seed[2422],seed[1157],seed[2818],seed[3369],seed[3188],seed[3212],seed[1936],seed[743],seed[779],seed[665],seed[2621],seed[3906],seed[657],seed[860],seed[306],seed[112],seed[1729],seed[774],seed[1535],seed[1387],seed[910],seed[2076],seed[2250],seed[413],seed[843],seed[1368],seed[1024],seed[1591],seed[4038],seed[2131],seed[2676],seed[1318],seed[1576],seed[854],seed[3456],seed[1838],seed[2239],seed[3177],seed[3652],seed[2154],seed[1983],seed[639],seed[111],seed[243],seed[629],seed[2273],seed[2300],seed[3321],seed[1691],seed[12],seed[1909],seed[2812],seed[1886],seed[567],seed[1295],seed[350],seed[1586],seed[450],seed[3409],seed[1781],seed[3962],seed[4060],seed[2641],seed[2932],seed[1610],seed[4072],seed[2121],seed[1847],seed[283],seed[3038],seed[3630],seed[189],seed[797],seed[3675],seed[133],seed[1526],seed[2595],seed[1094],seed[2845],seed[2808],seed[1661],seed[2433],seed[2775],seed[648],seed[2703],seed[1638],seed[527],seed[3446],seed[3545],seed[1429],seed[2788],seed[638],seed[3106],seed[1954],seed[898],seed[70],seed[1981],seed[2584],seed[3838],seed[2047],seed[2876],seed[3491],seed[3593],seed[706],seed[18],seed[1210],seed[3954],seed[1427],seed[127],seed[3951],seed[1672],seed[691],seed[749],seed[572],seed[4034],seed[3056],seed[2826],seed[813],seed[1099],seed[1302],seed[249],seed[2384],seed[1064],seed[3362],seed[2918],seed[1809],seed[2326],seed[1645],seed[4088],seed[2078],seed[179],seed[1650],seed[3883],seed[1864],seed[1912],seed[3975],seed[331],seed[109],seed[3173],seed[3257],seed[1021],seed[1456],seed[733],seed[3164],seed[3728],seed[2236],seed[653],seed[2288],seed[2188],seed[2416],seed[1989],seed[3952],seed[836],seed[3587],seed[2534],seed[1826],seed[2254],seed[613],seed[1702],seed[253],seed[120],seed[1979],seed[1760],seed[2564],seed[2637],seed[1160],seed[2900],seed[964],seed[1608],seed[3550],seed[2446],seed[3595],seed[4089],seed[562],seed[3122],seed[3907],seed[186],seed[3285],seed[3015],seed[3070],seed[1491],seed[292],seed[1153],seed[1609],seed[3093],seed[2152],seed[1643],seed[3104],seed[281],seed[40],seed[3941],seed[3606],seed[2752],seed[1335],seed[2803],seed[3688],seed[3897],seed[799],seed[3902],seed[3278],seed[4025],seed[2815],seed[468],seed[1209],seed[2533],seed[1622],seed[215],seed[2605],seed[583],seed[902],seed[1915],seed[1176],seed[1962],seed[1323],seed[2082],seed[3507],seed[859],seed[2695],seed[1304],seed[857],seed[905],seed[3225],seed[2160],seed[1816],seed[1402],seed[472],seed[823],seed[524],seed[2447],seed[3752],seed[980],seed[602],seed[3344],seed[3372],seed[2795],seed[3803],seed[1338],seed[4069],seed[982],seed[251],seed[2869],seed[1765],seed[2650],seed[3694],seed[427],seed[1253],seed[152],seed[3812],seed[1722],seed[3108],seed[1520],seed[311],seed[2569],seed[529],seed[977],seed[3025],seed[1592],seed[636],seed[2180],seed[3232],seed[293],seed[4044],seed[1628],seed[103],seed[1437],seed[3139],seed[2913],seed[2278],seed[2280],seed[3190],seed[875],seed[2111],seed[2714],seed[3567],seed[630],seed[3776],seed[246],seed[1399],seed[3939],seed[4056],seed[1107],seed[556],seed[1453],seed[3672],seed[1517],seed[2243],seed[336],seed[2935],seed[3319],seed[1935],seed[395],seed[2616],seed[3835],seed[1739],seed[3141],seed[1228],seed[563],seed[3283],seed[53],seed[2770],seed[3524],seed[201],seed[57],seed[3660],seed[948],seed[2353],seed[2041],seed[3631],seed[2130],seed[2436],seed[399],seed[1632],seed[2169],seed[280],seed[752],seed[3874],seed[3614],seed[1405],seed[320],seed[2158],seed[145],seed[976],seed[712],seed[1762],seed[3748],seed[1458],seed[2991],seed[2933],seed[3067],seed[3860],seed[1991],seed[2125],seed[1089],seed[3522],seed[3820],seed[2065],seed[36],seed[3789],seed[867],seed[2045],seed[3625],seed[695],seed[1286],seed[2875],seed[1311],seed[698],seed[1529],seed[545],seed[1128],seed[3352],seed[1795],seed[763],seed[116],seed[827],seed[3430],seed[3517],seed[1867],seed[2678],seed[619],seed[3990],seed[999],seed[3185],seed[1412],seed[3417],seed[349],seed[2837],seed[1140],seed[341],seed[3949],seed[2427],seed[3683],seed[50],seed[3144],seed[1310],seed[28],seed[943],seed[2014],seed[3486],seed[892],seed[528],seed[1103],seed[3731],seed[3687],seed[2940],seed[4039],seed[1792],seed[3199],seed[3037],seed[2066],seed[1705],seed[3716],seed[2186],seed[2660],seed[3733],seed[1197],seed[2166],seed[1756],seed[3147],seed[584],seed[1922],seed[2026],seed[3667],seed[1689],seed[2614],seed[3099],seed[1680],seed[49],seed[3588],seed[1759],seed[3821],seed[1439],seed[3057],seed[3330],seed[3131],seed[2737],seed[3503],seed[2997],seed[1347],seed[3314],seed[314],seed[2208],seed[808],seed[1334],seed[1397],seed[3244],seed[1046],seed[500],seed[347],seed[1395],seed[345],seed[1137],seed[3632],seed[2029],seed[371],seed[3339],seed[1240],seed[2490],seed[1623],seed[433],seed[946],seed[3485],seed[1613],seed[392],seed[734],seed[1504],seed[2459],seed[3428],seed[2836],seed[3501],seed[3610],seed[2283],seed[479],seed[3682],seed[1641],seed[2526],seed[2017],seed[2064],seed[4036],seed[3398],seed[2970],seed[3833],seed[1627],seed[2799],seed[1275],seed[3868],seed[304],seed[3434],seed[1278],seed[1279],seed[3348],seed[3512],seed[1522],seed[1749],seed[82],seed[128],seed[3925],seed[3754],seed[929],seed[3980],seed[610],seed[198],seed[1148],seed[1432],seed[2760],seed[2736],seed[969],seed[3496],seed[1919],seed[222],seed[1925],seed[671],seed[2322],seed[418],seed[1357],seed[1553],seed[2256],seed[3324],seed[1300],seed[2484],seed[3247],seed[2746],seed[965],seed[769],seed[2081],seed[1414],seed[1570],seed[1600],seed[2398],seed[3735],seed[1955],seed[4055],seed[3095],seed[1891],seed[2117],seed[512],seed[2864],seed[3197],seed[2059],seed[2221],seed[3921],seed[505],seed[660],seed[1150],seed[4028],seed[192],seed[2839],seed[1670],seed[2509],seed[2898],seed[782],seed[3917],seed[3575],seed[2723],seed[2697],seed[3686],seed[1236],seed[3499],seed[1665],seed[1818],seed[14],seed[2248],seed[3461],seed[1030],seed[3602],seed[2834],seed[3184],seed[259],seed[4012],seed[1131],seed[3282],seed[3965],seed[3742],seed[693],seed[2318],seed[2773],seed[3079],seed[742],seed[221],seed[3206],seed[3872],seed[459],seed[2073],seed[881],seed[2055],seed[380],seed[31],seed[3251],seed[662],seed[3351],seed[3546],seed[805],seed[338],seed[1988],seed[441],seed[1658],seed[791],seed[0],seed[137],seed[1621],seed[560],seed[1114],seed[3011],seed[4051],seed[503],seed[1440],seed[3198],seed[1224],seed[3101],seed[2444],seed[305],seed[1101],seed[1692],seed[815],seed[3645],seed[3696],seed[184],seed[144],seed[2167],seed[1519],seed[2645],seed[3890],seed[3695],seed[3354],seed[3691],seed[2168],seed[2448],seed[3730],seed[3120],seed[3214],seed[1679],seed[3679],seed[2912],seed[3117],seed[907],seed[3412],seed[1882],seed[1356],seed[728],seed[1465],seed[3127],seed[2506],seed[387],seed[1034],seed[2077],seed[2261],seed[1459],seed[2607],seed[853],seed[3337],seed[2298],seed[3192],seed[2463],seed[825],seed[1353],seed[373],seed[2139],seed[2822],seed[3663],seed[1582],seed[183],seed[839],seed[2343],seed[1596],seed[2562],seed[3829],seed[3787],seed[257],seed[2179],seed[3294],seed[2266],seed[2531],seed[3594],seed[3451],seed[844],seed[2783],seed[3792],seed[3992],seed[1798],seed[2833],seed[429],seed[802],seed[1196],seed[188],seed[3920],seed[2311],seed[1797],seed[784],seed[985],seed[3051],seed[9],seed[129],seed[44],seed[1175],seed[2395],seed[69],seed[2219],seed[3904],seed[1799],seed[3218],seed[1085],seed[796],seed[828],seed[1690],seed[118],seed[2787],seed[1676],seed[1881],seed[181],seed[1646],seed[2655],seed[158],seed[2916],seed[2625],seed[3227],seed[3670],seed[1256],seed[3304],seed[3073],seed[166],seed[3571],seed[3264],seed[3256],seed[2690],seed[3714],seed[1449],seed[2380],seed[2608],seed[456],seed[2052],seed[2781],seed[454],seed[272],seed[1289],seed[291],seed[901],seed[3378],seed[3222],seed[2434],seed[2975],seed[2917],seed[3072],seed[962],seed[756],seed[3857],seed[515],seed[3361],seed[1727],seed[3426],seed[1321],seed[3196],seed[2031],seed[3573],seed[1487],seed[1267],seed[2810],seed[3143],seed[1617],seed[2735],seed[212],seed[3438],seed[2780],seed[67],seed[1438],seed[3287],seed[2259],seed[3137],seed[235],seed[3750],seed[1277],seed[1259],seed[2209],seed[2282],seed[3740],seed[581],seed[2871],seed[3183],seed[2617],seed[2520],seed[2128],seed[1127],seed[2499],seed[2216],seed[3822],seed[2418],seed[1095],seed[2],seed[3521],seed[2230],seed[2303],seed[344],seed[3599],seed[4017],seed[3697],seed[2994],seed[3718],seed[1927],seed[1325],seed[3978],seed[861],seed[1163],seed[2681],seed[3246],seed[1180],seed[2659],seed[2571],seed[3404],seed[2269],seed[963],seed[1802],seed[1392],seed[3858],seed[475],seed[1416],seed[1514],seed[740],seed[2959],seed[924],seed[1467],seed[3163],seed[2575],seed[224],seed[1362],seed[504],seed[2794],seed[2604],seed[3782],seed[1785],seed[232],seed[1184],seed[2813],seed[1265],seed[606],seed[4029],seed[403],seed[709],seed[3995],seed[1179],seed[3841],seed[439],seed[2570],seed[2558],seed[3544],seed[838],seed[209],seed[485],seed[1067],seed[1044],seed[1580],seed[1173],seed[1447],seed[3930],seed[3458],seed[1743],seed[918],seed[3482],seed[1499],seed[470],seed[3813],seed[1464],seed[2613],seed[2241],seed[1488],seed[1862],seed[1483],seed[219],seed[2583],seed[1367],seed[3112],seed[1037],seed[353],seed[2831],seed[4006],seed[2858],seed[2175],seed[1509],seed[352],seed[2195],seed[3526],seed[1616],seed[1396],seed[2937],seed[759],seed[1768],seed[240],seed[1100],seed[1551],seed[2860],seed[3725],seed[2357],seed[2027],seed[3909],seed[2290],seed[1307],seed[3415],seed[780],seed[2973],seed[1742],seed[1369],seed[1328],seed[775],seed[758],seed[2423],seed[2734],seed[2574],seed[3064],seed[3910],seed[3474],seed[1857],seed[2846],seed[2715],seed[4094],seed[2372],seed[3489],seed[1109],seed[226],seed[2354],seed[1833],seed[480],seed[227],seed[921],seed[309],seed[2744],seed[787],seed[1422],seed[410],seed[2612],seed[1301],seed[1996],seed[3274],seed[522],seed[3692],seed[3425],seed[1455],seed[1376],seed[2748],seed[33],seed[1139],seed[3024],seed[1492],seed[329],seed[231],seed[3468],seed[1266],seed[711],seed[1250],seed[930],seed[1984],seed[1381],seed[2996],seed[444],seed[3018],seed[3266],seed[2670],seed[587],seed[490],seed[3242],seed[2624],seed[2927],seed[645],seed[2363],seed[1187],seed[4026],seed[754],seed[3781],seed[2165],seed[991],seed[2205],seed[2609],seed[2950],seed[3275],seed[1914],seed[492],seed[1855],seed[3288],seed[1612],seed[661],seed[3542],seed[2386],seed[396],seed[3449],seed[3086],seed[1726],seed[1326],seed[3862],seed[2319],seed[316],seed[4079],seed[550],seed[87],seed[3158],seed[837],seed[1027],seed[3250],seed[2701],seed[2331],seed[187],seed[2244],seed[2656],seed[4087],seed[2694],seed[3230],seed[3745],seed[1571],seed[3423],seed[1640],seed[1585],seed[2778],seed[1388],seed[1642],seed[1629],seed[1928],seed[230],seed[3179],seed[3662],seed[1308],seed[1566],seed[3578],seed[3026],seed[1965],seed[2896],seed[3793],seed[767],seed[2226],seed[1734],seed[2299],seed[3171],seed[2159],seed[1754],seed[2537],seed[2381],seed[981],seed[2136],seed[3472],seed[342],seed[2911],seed[1777],seed[2566],seed[1003],seed[579],seed[631],seed[13],seed[3320],seed[1892],seed[1997],seed[3062],seed[3012],seed[2477],seed[2848],seed[2590],seed[2338],seed[3736],seed[2197],seed[3926],seed[2840],seed[151],seed[2661],seed[3201],seed[2716],seed[3323],seed[2092],seed[30],seed[870],seed[3302],seed[1693],seed[1516],seed[1796],seed[3186],seed[3316],seed[156],seed[1410],seed[1012],seed[3429],seed[202],seed[689],seed[1283],seed[3867],seed[2116],seed[841],seed[2529],seed[612],seed[3022],seed[1011],seed[3987],seed[1557],seed[2948],seed[2790],seed[1126],seed[1942],seed[1306],seed[2265],seed[591],seed[2007],seed[3997],seed[2706],seed[620],seed[2974],seed[564],seed[1312],seed[3142],seed[1195],seed[3654],seed[2630],seed[2036],seed[2494],seed[294],seed[499],seed[2545],seed[2150],seed[1843],seed[3515],seed[1485],seed[2191],seed[2915],seed[2471],seed[2954],seed[3600],seed[3809],seed[961],seed[163],seed[1254],seed[3843],seed[1539],seed[2942],seed[940],seed[1827],seed[96],seed[1025],seed[3871],seed[1226],seed[3895],seed[140],seed[3033],seed[2192],seed[3153],seed[1595],seed[866],seed[1201],seed[3647],seed[3125],seed[3063],seed[3149],seed[1589],seed[2443],seed[2786],seed[481],seed[401],seed[1418],seed[3893],seed[3495],seed[3936],seed[1852],seed[3165],seed[594],seed[416],seed[3615],seed[1717],seed[3050],seed[1911],seed[2341],seed[2741],seed[2144],seed[2161],seed[3295],seed[2765],seed[738],seed[1830],seed[3948],seed[2025],seed[1682],seed[3381],seed[2011],seed[2776],seed[3601],seed[3306],seed[3769],seed[2667],seed[2049],seed[3296],seed[1206],seed[1398],seed[1811],seed[1384],seed[1663],seed[2749],seed[1877],seed[862],seed[2473],seed[2960],seed[2060],seed[973],seed[1614],seed[2557],seed[1272],seed[846],seed[1512],seed[781],seed[2342],seed[3336],seed[4027],seed[258],seed[2229],seed[2387],seed[1169],seed[1124],seed[2989],seed[3317],seed[748],seed[1460],seed[2669],seed[2435],seed[2816],seed[148],seed[3152],seed[3702],seed[1967],seed[2987],seed[960],seed[3475],seed[607],seed[2222],seed[2925],seed[2789],seed[108],seed[1834],seed[3582],seed[2591],seed[3268],seed[1339],seed[351],seed[3592],seed[1309],seed[1284],seed[959],seed[3175],seed[3031],seed[3847],seed[732],seed[2718],seed[3393],seed[1500],seed[4037],seed[3574],seed[2393],seed[3457],seed[2126],seed[2437],seed[2142],seed[2048],seed[372],seed[2091],seed[3366],seed[1031],seed[3103],seed[3454],seed[2177],seed[549],seed[2618],seed[3918],seed[1288],seed[1270],seed[35],seed[967],seed[1652],seed[2333],seed[3756],seed[2348],seed[3309],seed[2185],seed[664],seed[2992],seed[883],seed[1649],seed[3328],seed[900],seed[2072],seed[1771],seed[2184],seed[3642],seed[1587],seed[2213],seed[1873],seed[865],seed[2367],seed[1974],seed[2420],seed[1869],seed[2983],seed[1141],seed[3035],seed[3200],seed[1933],seed[3333],seed[2441],seed[697],seed[1022],seed[2492],seed[1712],seed[2895],seed[3097],seed[2504],seed[2881],seed[674],seed[223],seed[771],seed[2668],seed[3559],seed[1461],seed[2401],seed[713],seed[950],seed[3280],seed[1822],seed[1916],seed[464],seed[2689],seed[4008],seed[3796],seed[1042],seed[1448],seed[3480],seed[1161],seed[414],seed[75],seed[2792],seed[3887],seed[1704],seed[538],seed[3135],seed[92],seed[3611],seed[708],seed[303],seed[1494],seed[3493],seed[58],seed[2408],seed[2552],seed[393],seed[1002],seed[3347],seed[317],seed[2083],seed[2643],seed[3802],seed[3580],seed[2346],seed[1956],seed[1247],seed[3410],seed[1041],seed[3224],seed[2249],seed[2796],seed[1386],seed[995],seed[1478],seed[3661],seed[3955],seed[2947],seed[1923],seed[3643],seed[2855],seed[1181],seed[2811],seed[2798],seed[1725],seed[2977],seed[2090],seed[1102],seed[745],seed[2050],seed[1212],seed[2633],seed[3659],seed[2934],seed[2138],seed[3374],seed[168],seed[3481],seed[1377],seed[904],seed[375],seed[3986],seed[2622],seed[1049],seed[3523],seed[1066],seed[1724],seed[714],seed[1975],seed[3094],seed[2511],seed[2536],seed[457],seed[3259],seed[2291],seed[1213],seed[2647],seed[634],seed[534],seed[3300],seed[1669],seed[795],seed[3514],seed[274],seed[3689],seed[822],seed[1874],seed[1078],seed[210],seed[2003],seed[290],seed[104],seed[376],seed[1020],seed[3401],seed[2698],seed[234],seed[1394],seed[16],seed[390],seed[1477],seed[1987],seed[287],seed[3484],seed[3039],seed[2432],seed[269],seed[942],seed[816],seed[3356],seed[3519],seed[3435],seed[2198],seed[2677],seed[102],seed[1502],seed[1428],seed[2733],seed[1907],seed[2593],seed[2057],seed[3773],seed[86],seed[2100],seed[736],seed[3828],seed[1808],seed[869],seed[1409],seed[3174],seed[2033],seed[2666],seed[1331],seed[3861],seed[3014],seed[1720],seed[3036],seed[176],seed[1425],seed[3360],seed[3269],seed[2938],seed[313],seed[3045],seed[1884],seed[1906],seed[2874],seed[2068],seed[729],seed[3145],seed[2555],seed[2356],seed[886],seed[2133],seed[2944],seed[2337],seed[1993],seed[2865],seed[3617],seed[1647],seed[3439],seed[2493],seed[3864],seed[1770],seed[1684],seed[2360],seed[4033],seed[2646],seed[997],seed[725],seed[237],seed[1863],seed[164],seed[3450],seed[673],seed[25],seed[1593],seed[2464],seed[1918],seed[1681],seed[3935],seed[3923],seed[2628],seed[2549],seed[817],seed[642],seed[465],seed[161],seed[65],seed[3786],seed[2971],seed[2686],seed[2301],seed[2887],seed[333],seed[700],seed[3896],seed[278],seed[1424],seed[2882],seed[1872],seed[1934],seed[2867],seed[1594],seed[3138],seed[3349],seed[3263],seed[718],seed[2129],seed[2215],seed[1578],seed[3898],seed[3364],seed[1075],seed[531],seed[2528],seed[141],seed[1769],seed[383],seed[2252],seed[4068],seed[2482],seed[2019],seed[1940],seed[1832],seed[3541],seed[3946],seed[1010],seed[1950],seed[677],seed[1687],seed[453],seed[3297],seed[340],seed[43],seed[3963],seed[2147],seed[1207],seed[355],seed[1673],seed[2654],seed[3189],seed[3416],seed[1220],seed[1352],seed[2606],seed[2964],seed[3020],seed[1382],seed[1451],seed[3237],seed[3226],seed[3272],seed[2885],seed[2094],seed[134],seed[770],seed[2231],seed[1084],seed[2276],seed[1791],seed[3953],seed[4000],seed[3966],seed[4065],seed[312],seed[2560],seed[248],seed[2889],seed[2310],seed[3815],seed[2980],seed[1055],seed[3508],seed[3299],seed[565],seed[3403],seed[3973],seed[3502],seed[3167],seed[2635],seed[3466],seed[357],seed[3156],seed[296],seed[1846],seed[1840],seed[1132],seed[2819],seed[3612],seed[95],seed[2012],seed[1182],seed[452],seed[1958],seed[100],seed[628],seed[2768],seed[1930],seed[3950],seed[2611],seed[2649],seed[54],seed[2951],seed[3445],seed[1350],seed[510],seed[1198],seed[3724],seed[3794],seed[2880],seed[88],seed[894],seed[1482],seed[1948],seed[1801],seed[702],seed[8],seed[451],seed[2472],seed[2204],seed[692],seed[1960],seed[2945],seed[2268],seed[2228],seed[2620],seed[954],seed[1230],seed[2430],seed[4024],seed[81],seed[588],seed[2227],seed[319],seed[1341],seed[2801],seed[107],seed[1546],seed[1775],seed[1949],seed[658],seed[3157],seed[2350],seed[359],seed[966],seed[3010],seed[245],seed[4059],seed[1992],seed[2108],seed[1573],seed[3510],seed[3389],seed[1841],seed[2523],seed[2114],seed[277],seed[2355],seed[2009],seed[1708],seed[3982],seed[2097],seed[297],seed[914],seed[2894],seed[831],seed[2502],seed[22],seed[97],seed[3098],seed[1471],seed[2352],seed[2086],seed[2955],seed[1233],seed[3365],seed[150],seed[2651],seed[3525],seed[2827],seed[2598],seed[1147],seed[3974],seed[1199],seed[126],seed[3607],seed[3028],seed[1943],seed[2307],seed[1237],seed[3551],seed[1985],seed[1285],seed[182],seed[2403],seed[1214],seed[3845],seed[4092],seed[250],seed[204],seed[2705],seed[1462],seed[3312],seed[2485],seed[2619],seed[3915],seed[1543],seed[1696],seed[647],seed[876],seed[2178],seed[878],seed[366],seed[3999],seed[604],seed[1071],seed[3058],seed[3819],seed[3081],seed[2292],seed[1966],seed[1457],seed[268],seed[2862],seed[2253],seed[580],seed[1844],seed[2683],seed[3598],seed[2340],seed[2998],seed[2242],seed[1648],seed[672],seed[467],seed[3699],seed[1361],seed[1446],seed[3676],seed[2389],seed[1229],seed[3554],seed[3181],seed[3091],seed[3622],seed[3996],seed[2685],seed[788],seed[2507],seed[46],seed[2449],seed[2406],seed[3215],seed[3436],seed[3100],seed[2892],seed[2627],seed[3068],seed[2370],seed[3009],seed[1837],seed[798],seed[2747],seed[3649],seed[2487],seed[1166],seed[398],seed[2731],seed[1978],seed[2275],seed[1401],seed[1655],seed[3236],seed[1825],seed[2196],seed[3976],seed[3041],seed[1496],seed[2551],seed[2272],seed[2383],seed[3090],seed[933],seed[2853],seed[1659],seed[2417],seed[1990],seed[949],seed[270],seed[1611],seed[1635],seed[1372],seed[2601],seed[2402],seed[2724],seed[688],seed[701],seed[814],seed[346],seed[737],seed[3194],seed[2379],seed[1366],seed[1639],seed[1243],seed[2720],seed[680],seed[3658],seed[94],seed[415],seed[2738],seed[1],seed[2688],seed[998],seed[59],seed[2118],seed[986],seed[1248],seed[576],seed[1186],seed[2211],seed[927],seed[3140],seed[1730],seed[2388],seed[739],seed[3082],seed[1231],seed[1653],seed[1081],seed[1105],seed[2329],seed[2907],seed[513],seed[703],seed[1346],seed[3712],seed[1490],seed[557],seed[1737],seed[4022],seed[2691],seed[852],seed[241],seed[2458],seed[2514],seed[1565],seed[2409],seed[2772],seed[1503],seed[3807],seed[2730],seed[2993],seed[1913],seed[2232],seed[2638],seed[945],seed[1773],seed[3539],seed[721],seed[4042],seed[497],seed[2442],seed[3931],seed[2847],seed[3869],seed[365],seed[207],seed[443],seed[821],seed[3397],seed[3770],seed[2106],seed[3407],seed[1820],seed[2439],seed[426],seed[877],seed[3693],seed[1445],seed[682],seed[936],seed[1794],seed[3804],seed[1783],seed[1929],seed[1219],seed[256],seed[3556],seed[2465],seed[681],seed[2956],seed[3238],seed[1544],seed[4003],seed[3638],seed[548],seed[3518],seed[3487],seed[1941],seed[696],seed[2234],seed[2728],seed[411],seed[1545],seed[388],seed[3881],seed[1466],seed[1851],seed[430],seed[167],seed[1061],seed[3],seed[3327],seed[1698],seed[3281],seed[3771],seed[820],seed[21],seed[1480],seed[327],seed[2692],seed[279],seed[2759],seed[1697],seed[2902],seed[1633],seed[521],seed[89],seed[3772],seed[3455],seed[1555],seed[496],seed[3814],seed[3856],seed[449],seed[404],seed[2967],seed[1938],seed[84],seed[3678],seed[2854],seed[85],seed[1415],seed[508],seed[1953],seed[73],seed[142],seed[715],seed[3110],seed[1603],seed[1814],seed[4086],seed[2115],seed[807],seed[2893],seed[911],seed[1865],seed[753],seed[3880],seed[1531],seed[750],seed[1106],seed[3540],seed[76],seed[1959],seed[91],seed[3816],seed[2093],seed[1900],seed[3205],seed[726],seed[934],seed[2016],seed[4058],seed[578],seed[1878],seed[3870],seed[1527],seed[3913],seed[2722],seed[2756],seed[56],seed[4067],seed[2258],seed[147],seed[3380],seed[3779],seed[405],seed[2704],seed[1699],seed[2190],seed[2371],seed[2022],seed[298],seed[2580],seed[3055],seed[1167],seed[2217],seed[3359],seed[328],seed[3969],seed[1508],seed[1706],seed[970],seed[4047],seed[1257],seed[60],seed[381],seed[1518],seed[3007],seed[1009],seed[3768],seed[4073],seed[4045],seed[3467],seed[1108],seed[507],seed[2755],seed[3129],seed[3561],seed[3985],seed[3746],seed[1533],seed[125],seed[3788],seed[667],seed[2286],seed[3853],seed[1736],seed[4070],seed[1174],seed[2453],seed[2474],seed[2921],seed[2260],seed[2067],seed[3379],seed[3154],seed[1964],seed[4048],seed[2470],seed[2366],seed[551],seed[2431],seed[2039],seed[3029],seed[3160],seed[1764],seed[3303],seed[1324],seed[2173],seed[1242],seed[2143],seed[1537],seed[3326],seed[3030],seed[2376],seed[2425],seed[423],seed[3270],seed[1719],seed[3938],seed[1607],seed[539],seed[2302],seed[1619],seed[3075],seed[707],seed[951],seed[2708],seed[618],seed[420],seed[2235],seed[2120],seed[1731],seed[3452],seed[2270],seed[1876],seed[1400],seed[3161],seed[735],seed[1217],seed[979],seed[2127],seed[3916],seed[362],seed[42],seed[1750],seed[2626],seed[1728],seed[1098],seed[2554],seed[2824],seed[3671],seed[2438],seed[3343],seed[773],seed[1403],seed[1858],seed[3558],seed[3836],seed[1282],seed[2214],seed[2218],seed[1436],seed[746],seed[1744],seed[675],seed[1097],seed[29],seed[3584],seed[228],seed[2962],seed[473],seed[1893],seed[1807],seed[760],seed[310],seed[616],seed[3644],seed[121],seed[623],seed[1470],seed[2028],seed[238],seed[1569],seed[3402],seed[407],seed[3492],seed[832],seed[2579],seed[4095],seed[3229],seed[4019],seed[1572],seed[683],seed[3276],seed[1407],seed[2856],seed[590],seed[1281],seed[247],seed[3054],seed[793],seed[27],seed[3134],seed[2396],seed[872],seed[649],seed[1315],seed[2600],seed[932],seed[903],seed[200],seed[2986],seed[3763],seed[2002],seed[3989],seed[2957],seed[1146],seed[1391],seed[3052],seed[3945],seed[2984],seed[1019],seed[687],seed[3709],seed[1417],seed[3624],seed[1047],seed[2546],seed[3826],seed[1441],seed[254],seed[3074],seed[1803],seed[2508],seed[2156],seed[2674],seed[445],seed[1070],seed[178],seed[442],seed[2515],seed[1969],seed[7],seed[1711],seed[422],seed[2246],seed[543],seed[694],seed[428],seed[3548],seed[2561],seed[2483],seed[367],seed[1709],seed[2004],seed[3797],seed[1973],seed[1524],seed[2979],seed[19],seed[199],seed[1303],seed[3879],seed[2978],seed[2255],seed[2793],seed[923],seed[1761],seed[2965],seed[3665],seed[3208],seed[3784],seed[197],seed[3498],seed[379],seed[1443],seed[4057],seed[1133],seed[2308],seed[4085],seed[1618],seed[3531],seed[1668],seed[3605],seed[2632],seed[978],seed[2936],seed[195],seed[3078],seed[1261],seed[2563],seed[1757],seed[1856],seed[840],seed[2577],seed[863],seed[1050],seed[3597],seed[1129],seed[2053],seed[3527],seed[2582],seed[51],seed[3533],seed[2553],seed[3706],seed[3080],seed[1547],seed[1921],seed[3119],seed[261],seed[3656],seed[690],seed[2061],seed[3395],seed[421],seed[3210],seed[540],seed[3774],seed[1980],seed[2105],seed[1378],seed[1143],seed[812],seed[3008],seed[3353],seed[678],seed[3405],seed[1297],seed[2141],seed[2547],seed[2804],seed[2365],seed[2929],seed[1784],seed[1280],seed[3855],seed[2399],seed[1534],seed[1790],seed[2101],seed[656],seed[585],seed[1605],seed[307],seed[322],seed[1014],seed[764],seed[2194],seed[1238],seed[2405],seed[596],seed[3576],seed[3943],seed[1707],seed[171],seed[2306],seed[2132],seed[286],seed[890],seed[3705],seed[3187],seed[3717],seed[384],seed[855],seed[1332],seed[130],seed[1013],seed[1389],seed[52],seed[2429],seed[493],seed[3979],seed[974],seed[3875],seed[3396],seed[1821],seed[3209],seed[633],seed[177],seed[2394],seed[3673],seed[321],seed[3604],seed[3291],seed[1245],seed[893],seed[4035],seed[3536],seed[3345],seed[2522],seed[611],seed[3957],seed[858],seed[2368],seed[1671],seed[1848],seed[1435],seed[2807],seed[1336],seed[2295],seed[1040],seed[397],seed[3873],seed[3202],seed[1191],seed[446],seed[2878],seed[2629],seed[1880],seed[1342],seed[4050],seed[1134],seed[2153],seed[236],seed[2671],seed[3901],seed[3719],seed[1894],seed[2713],seed[2914],seed[2615],seed[3831],seed[3703],seed[2518],seed[553],seed[1452],seed[218],seed[761],seed[983],seed[2838],seed[3087],seed[2001],seed[193],seed[654],seed[3775],seed[3207],seed[1778],seed[285],seed[339],seed[888],seed[1898],seed[3783],seed[3749],seed[3560],seed[1234],seed[2032],seed[2358],seed[1902],seed[1255],seed[1804],seed[2931],seed[2763],seed[830],seed[3377],seed[2411],seed[162],seed[3669],seed[1365],seed[2334],seed[1379],seed[3690],seed[23],seed[988],seed[334],seed[233],seed[3555],seed[3633],seed[2919],seed[2410],seed[3422],seed[2155],seed[3476],seed[3981],seed[2901],seed[48],seed[3668],seed[3367],seed[644],seed[356],seed[2870],seed[2538],seed[1637],seed[776],seed[3228],seed[1971],seed[2104],seed[1317],seed[1004],seed[3811],seed[1944],seed[3998],seed[3292],seed[1138],seed[1287],seed[2099],seed[3385],seed[2098],seed[139],seed[364],seed[2021],seed[1530],seed[1497],seed[3727],seed[3721],seed[1168],seed[1244],seed[1130],seed[2725],seed[1758],seed[2985],seed[2585],seed[3453],seed[3892],seed[2263],seed[3136],seed[1866],seed[806],seed[2497],seed[315],seed[1029],seed[3859],seed[1112],seed[939],seed[3130],seed[1120],seed[2426],seed[3929],seed[1889],seed[1563],seed[913],seed[2884],seed[801],seed[3500],seed[1835],seed[1767],seed[785],seed[2825],seed[595],seed[3162],seed[778],seed[3967],seed[2700],seed[1154],seed[1232],seed[1812],seed[2392],seed[3248],seed[3830],seed[1986],seed[1091],seed[3350],seed[3168],seed[509],seed[3221],seed[2203],seed[2527],seed[3260],seed[532],seed[3220],seed[2440],seed[2843],seed[1561],seed[3027],seed[1532],seed[3239],seed[1904],seed[917],seed[850],seed[2930],seed[947],seed[386],seed[3707],seed[1205],seed[3739],seed[3105],seed[3844],seed[1806],seed[3817],seed[2806],seed[2247],seed[1273],seed[1235],seed[255],seed[824],seed[3085],seed[3651],seed[1276],seed[2897],seed[216],seed[3341],seed[1156],seed[4021],seed[3133],seed[463],seed[2008],seed[2293],seed[2468],seed[206],seed[1579],seed[818],seed[1732],seed[3443],seed[2530],seed[32],seed[3441],seed[1700],seed[915],seed[2777],seed[2135],seed[3933],seed[953],seed[1701],seed[3114],seed[498],seed[3790],seed[2495],seed[2206],seed[157],seed[598],seed[3919],seed[2193],seed[514],seed[165],seed[3734],seed[2157],seed[1223],seed[4023],seed[2817],seed[39],seed[3623],seed[2802],seed[3572],seed[1656],seed[3148],seed[2849],seed[1420],seed[3650],seed[3253],seed[271],seed[1718],seed[358],seed[1963],seed[3286],seed[1604],seed[931],seed[2567],seed[3069],seed[1149],seed[2037],seed[3908],seed[3937],seed[2412],seed[1860],seed[555],seed[4071],seed[2886],seed[2359],seed[1776],seed[2774],seed[3490],seed[1899],seed[2262],seed[1495],seed[3254],seed[3241],seed[1385],seed[2739],seed[2751],seed[1875],seed[2289],seed[502],seed[1871],seed[747],seed[3488],seed[2267],seed[3406],seed[768],seed[1738],seed[1525],seed[3764],seed[3808],seed[1296],seed[3700],seed[1774],seed[1828],seed[289],seed[1383],seed[1327],seed[64],seed[891],seed[78],seed[1716],seed[2102],seed[3370],seed[517],seed[1678],seed[2923],seed[3626],seed[755],seed[676],seed[1033],seed[6],seed[1360],seed[2320],seed[2279],seed[2754],seed[605],seed[2457],seed[2820],seed[2664],seed[3577],seed[3537],seed[2890],seed[484],seed[1513],seed[1017],seed[546],seed[447],seed[1782],seed[265],seed[10],seed[525],seed[717],seed[1789],seed[3191],seed[3528],seed[1810],seed[987],seed[2095],seed[4016],seed[2451],seed[3387],seed[2565],seed[4014],seed[845],seed[2764],seed[3761],seed[2148],seed[1599],seed[3427],seed[1686],seed[2220],seed[751],seed[3262],seed[1861],seed[1155],seed[2758],seed[1073],seed[3569],seed[3905],seed[11],seed[2044],seed[2103],seed[47],seed[864],seed[3180],seed[252],seed[2005],seed[264],seed[3128],seed[3338],seed[3219],seed[3096],seed[3373],seed[3960],seed[993],seed[2559],seed[2369],seed[2982],seed[3922],seed[3066],seed[1710],seed[180],seed[2062],seed[3799],seed[3780],seed[4020],seed[1079],seed[1111],seed[885],seed[1208],seed[1080],seed[2109],seed[3565],seed[93],seed[242],seed[3016],seed[1348],seed[3590],seed[3109],seed[3315],seed[1479],seed[3390],seed[2088],seed[3083],seed[3944],seed[518],seed[573],seed[436],seed[3657],seed[3408],seed[4049],seed[757],seed[632],seed[952],seed[3509],seed[1060],seed[45],seed[110],seed[3150],seed[4063],seed[834],seed[3603],seed[1145],seed[1069],seed[3471],seed[1688],seed[523],seed[3557],seed[811],seed[723],seed[2024],seed[804],seed[1897],seed[2336],seed[2785],seed[1982],seed[3653],seed[124],seed[1723],seed[3400],seed[955],seed[3641],seed[2397],seed[2578],seed[1746],seed[3115],seed[3852],seed[3267],seed[1552],seed[922],seed[3383],seed[136],seed[3616],seed[363],seed[3543],seed[3534],seed[3609],seed[205],seed[1116],seed[2377],seed[1588],seed[1703],seed[975],seed[3701],seed[2210],seed[2035],seed[2762],seed[1442],seed[1473],seed[3447],seed[2013],seed[1575],seed[2652],seed[2480],seed[1121],seed[719],seed[2709],seed[2966],seed[4061],seed[3988],seed[3755],seed[3293],seed[2257],seed[2390],seed[1188],seed[2866],seed[3504],seed[3233],seed[3332],seed[260],seed[2588],seed[3968],seed[1314],seed[3346],seed[2414],seed[2682],seed[488],seed[458],seed[3203],seed[1952],seed[2469],seed[400],seed[637],seed[3310],seed[1463],seed[906],seed[66],seed[2317],seed[494],seed[3621],seed[849],seed[2910],seed[874],seed[727],seed[1606],seed[643],seed[434],seed[668],seed[3704],seed[2673],seed[2112],seed[2501],seed[1651],seed[2745],seed[1074],seed[3563],seed[1337],seed[374],seed[3713],seed[1831],seed[552],seed[3851],seed[1344],seed[3047],seed[2074],seed[1558],seed[1426],seed[3664],seed[1135],seed[2767],seed[1051],seed[1117],seed[3318],seed[1164],seed[330],seed[1489],seed[220],seed[651],seed[1215],seed[1577],seed[406],seed[3473],seed[2455],seed[2475],seed[1032],seed[762],seed[3766],seed[3170],seed[882],seed[324],seed[1125],seed[1511],seed[2750],seed[3411],seed[2122],seed[4030],seed[1358],seed[2452],seed[3903],seed[2510],seed[2850],seed[1076],seed[1045],seed[2535],seed[2642],seed[2640],seed[1054],seed[24],seed[1419],seed[1824],seed[2233],seed[972],seed[99],seed[1330],seed[3738],seed[2539],seed[1674],seed[1354],seed[437],seed[2707],seed[2344],seed[2328],seed[990],seed[1528],seed[2597],seed[38],seed[1747],seed[3715],seed[1292],seed[2648],seed[2503],seed[3759],seed[1088],seed[2592],seed[2189],seed[1193],seed[2174],seed[1241],seed[1486],seed[3970],seed[3023],seed[2952],seed[318],seed[868],seed[2586],seed[1829],seed[4053],seed[1839],seed[3371],seed[2237],seed[394],seed[1252],seed[1068],seed[716],seed[213],seed[1677],seed[3494],seed[1849],seed[1026],seed[3102],seed[3795],seed[1926],seed[956],seed[3666],seed[3591],seed[1995],seed[2085],seed[1375],seed[2345],seed[2466],seed[2162],seed[3866],seed[79],seed[1931],seed[2711],seed[2672],seed[3325],seed[2809],seed[586],seed[2873],seed[2137],seed[2525],seed[2324],seed[1917],seed[2069],seed[2456],seed[2314],seed[1890],seed[3618],seed[3092],seed[368],seed[1316],seed[650],seed[614],seed[2313],seed[2224],seed[1968],seed[469],seed[1190],seed[3640],seed[1887],seed[3399],seed[1264],seed[2861],seed[627],seed[670],seed[460],seed[1634],seed[2800],seed[2572],seed[1222],seed[2462],seed[1225],seed[2717],seed[941],seed[20],seed[2378],seed[3111],seed[3358],seed[2602],seed[273],seed[1946],seed[1431],seed[3538],seed[2419],seed[1836],seed[377],seed[3848],seed[471],seed[3284],seed[2134],seed[570],seed[2023],seed[391],seed[3357],seed[3886],seed[448],seed[1110],seed[786],seed[2599],seed[2264],seed[626],seed[2251],seed[3947],seed[2928],seed[3322],seed[2335],seed[1178],seed[2883],seed[3639],seed[5],seed[3891],seed[879],seed[2187],seed[871],seed[1615],seed[535],seed[1355],seed[61],seed[1787],seed[2908],seed[772],seed[2176],seed[1505],seed[3386],seed[1421],seed[3088],seed[2784],seed[1521],seed[3927],seed[3235],seed[1484],seed[3155],seed[1299],seed[343],seed[1183],seed[3271],seed[2926],seed[2404],seed[2461],seed[1994],seed[3581],seed[2309],seed[2240],seed[615],seed[873],seed[2505],seed[2743],seed[1598],seed[2071],seed[3223],seed[4080],seed[3849],seed[474],seed[1654],seed[1883],seed[154],seed[3732],seed[1583],seed[155],seed[3674],seed[3424],seed[1083],seed[1434],seed[1721],seed[800],seed[1788],seed[378],seed[1903],seed[3777],seed[608],seed[1685],seed[1349],seed[1568],seed[2000],seed[3912],seed[3723],seed[2428],seed[3431],seed[169],seed[2587],seed[2467],seed[1077],seed[810],seed[1329],seed[2476],seed[2863],seed[1374],seed[3132],seed[803],seed[1657],seed[2823],seed[170],seed[1481],seed[1581],seed[369],seed[944],seed[2969],seed[686],seed[173],seed[2146],seed[2990],seed[3301],seed[710],seed[895],seed[2171],seed[4052],seed[1567],seed[3042],seed[114],seed[1028],seed[1239],seed[1062],seed[106],seed[4013],seed[2362],seed[71],seed[1444],seed[1268],seed[2662],seed[3469],seed[295],seed[1142],seed[574],seed[1056],seed[1177],seed[2968],seed[3991],seed[3720],seed[4076],seed[3568],seed[3977],seed[3737],seed[3758],seed[1104],seed[3884],seed[4064],seed[335],seed[288],seed[1507],seed[3388],seed[1320],seed[600],seed[1910],seed[2163],seed[2075],seed[1823],seed[2906],seed[3961],seed[994],seed[537],seed[1291],seed[3076],seed[3124],seed[2972],seed[466],seed[1113],seed[3307],seed[3846],seed[3801],seed[2481],seed[4007],seed[2145],seed[663],seed[2124],seed[3899],seed[3585],seed[1171],seed[3497],seed[501],seed[3553],seed[175],seed[3046],seed[666],seed[2544],seed[3255],seed[880],seed[3635],seed[3722],seed[3204],seed[2512],seed[1805],seed[3375],seed[3084],seed[2170],seed[3636],seed[4090],seed[2486],seed[2548],seed[3940],seed[1694],seed[3277],seed[3532],seed[2719],seed[601],seed[1772],seed[262],seed[3579],seed[1817],seed[2953],seed[3470],seed[1850],seed[519],seed[2323],seed[2151],seed[3854],seed[1072],seed[916],seed[2835],seed[3684],seed[4018],seed[3744],seed[1868],seed[2872],seed[1845],seed[1574],seed[2107],seed[3172],seed[2710],seed[3448],seed[3876],seed[1541],seed[4032],seed[3342],seed[1018],seed[3934],seed[989],seed[1048],seed[1905],seed[1118],seed[3984],seed[724],seed[2183],seed[3432],seed[113],seed[3619],seed[1560],seed[2821],seed[3460],seed[3298],seed[2277],seed[101],seed[3824],seed[3000],seed[3017],seed[3993],seed[1870],seed[3972],seed[2271],seed[3477],seed[4081],seed[1059],seed[2963],seed[2634],seed[847],seed[2687],seed[3392],seed[1998],seed[2415],seed[848],seed[1413],seed[2859],seed[3726],seed[2140],seed[1165],seed[483],seed[1813],seed[935],seed[2988],seed[4066],seed[143],seed[300],seed[1590],seed[3549],seed[2330],seed[1038],seed[1185],seed[2550],seed[589],seed[2769],seed[511],seed[4084],seed[856],seed[646],seed[2532],seed[3520],seed[1584],seed[3440],seed[2382],seed[3005],seed[1380],seed[1536],seed[105],seed[730],seed[896],seed[282],seed[1170],seed[2351],seed[1430],seed[3065],seed[2294],seed[1493],seed[3832],seed[432],seed[1472],seed[361],seed[1390],seed[731],seed[3040],seed[2779],seed[160],seed[2596],seed[2653],seed[83],seed[217],seed[2056],seed[655],seed[1675],seed[2888],seed[174],seed[2413],seed[3118],seed[1119],seed[641],seed[2844],seed[968],seed[1260],seed[3414],seed[370],seed[3583],seed[3878],seed[971],seed[558],seed[2500],seed[777],seed[4],seed[2832],seed[789],seed[2757],seed[2791],seed[3911],seed[1475],seed[3767],seed[766],seed[1468],seed[3680],seed[495],seed[263],seed[1957],seed[3620],seed[417],seed[1664],seed[3837],seed[1364],seed[2842],seed[1096],seed[835],seed[1052],seed[1246],seed[559],seed[3331],seed[122],seed[3478],seed[2516],seed[229],seed[1745],seed[2123],seed[489],seed[419],seed[4075],seed[2905],seed[765],seed[652],seed[2164],seed[2200],seed[3747],seed[1542],seed[2051],seed[3234],seed[897],seed[541],seed[1039],seed[2904],seed[214],seed[2297],seed[194],seed[2766],seed[3159],seed[2364],seed[2517],seed[3760],seed[3800],seed[1433],seed[3060],seed[2042],seed[15],seed[3071],seed[2899],seed[2321],seed[1158],seed[2038],seed[2521],seed[3289],seed[1498],seed[2287],seed[3547],seed[55],seed[3249],seed[1932],seed[3959],seed[2006],seed[1947],seed[1780],seed[3685],seed[2782],seed[3634],seed[2663],seed[3126],seed[2080],seed[3308],seed[3178],seed[2070],seed[3313],seed[302],seed[1227],seed[3827],seed[2828],seed[984],seed[705],seed[2096],seed[244],seed[919],seed[4002],seed[2084],seed[2316],seed[2922],seed[196],seed[3791],seed[2043],seed[547],seed[3513],seed[3608],seed[3290],seed[669],seed[3710],seed[2920],seed[462],seed[17],seed[3535],seed[3176],seed[1005],seed[299],seed[3279],seed[2496],seed[4078],seed[3741],seed[3211],seed[62],seed[1920],seed[912],seed[1660],seed[571],seed[1406],seed[4004],seed[1136],seed[1371],seed[131],seed[2498],seed[3646],seed[431],seed[3243],seed[2058],seed[1601],seed[1901],seed[926],seed[829],seed[4009],seed[2305],seed[2087],seed[3894],seed[958],seed[2540],seed[599],seed[1842],seed[3465],seed[925],seed[2868],seed[2644],seed[225],seed[2581],seed[440],seed[3698],seed[1819],seed[1293],seed[2304],seed[1800],seed[1854],seed[3169],seed[4082],seed[435],seed[3442],seed[98],seed[3419],seed[609],seed[533],seed[593],seed[1715],seed[1393],seed[568],seed[2631],seed[625],seed[908],seed[37],seed[149],seed[2753],seed[3273],seed[3340],seed[1087],seed[1262],seed[1298],seed[3433],seed[3677],seed[2238],seed[1370],seed[842],seed[2639],seed[3865],seed[577],seed[1786],seed[3382],seed[412],seed[275],seed[3505],seed[3900],seed[1501],seed[3265],seed[2407],seed[3413],seed[3363],seed[185],seed[1319],seed[1713],seed[3217],seed[2460],seed[3418],seed[2312],seed[3863],seed[520],seed[2202],seed[1007],seed[809],seed[3708],seed[3971],seed[478],seed[1620],seed[461],seed[3019],seed[575],seed[2841],seed[3765],seed[2015],seed[4001],seed[1469],seed[1015],seed[1151],seed[3810],seed[2675],seed[135],seed[2172],seed[2576],seed[337],seed[2761],seed[1093],seed[1753],seed[506],seed[1879],seed[3627],seed[530],seed[26],seed[138],seed[617],seed[3586],seed[1667],seed[3121],seed[1644],seed[90],seed[408],seed[3166],seed[3003],seed[3805],seed[3994],seed[1597],seed[4091],seed[2851],seed[3258],seed[1082],seed[1815],seed[1351],seed[2603],seed[2636],seed[2797],seed[1562],seed[1194],seed[2079],seed[635],seed[191],seed[2361],seed[622],seed[3355],seed[2721],seed[2696],seed[3061],seed[385],seed[889],seed[1008],seed[3942],seed[704],seed[2740],seed[2941],seed[3566],seed[2089],seed[1115],seed[2285],seed[621],seed[790],seed[516],seed[826],seed[792],seed[2729],seed[3564],seed[833],seed[3245],seed[2857],seed[1908],seed[2374],seed[2223],seed[3743],seed[1559],seed[3182],seed[2054],seed[3753],seed[1853],seed[1016],seed[1972],seed[2046],seed[1631],seed[2225],seed[1333],seed[3757],seed[3013],seed[424],seed[409],seed[1203],seed[1290],seed[1454],seed[2981],seed[2589],seed[2542],seed[2949],seed[1006],seed[1506],seed[3956],seed[1123],seed[3004],seed[1793],seed[34],seed[1666],seed[1204],seed[382],seed[1221],seed[2742],seed[1294],seed[3842],seed[2347],seed[3637],seed[3818],seed[624],seed[3762],seed[2010],seed[1554],seed[119],seed[2281],seed[323],seed[2829],seed[2877],seed[3479],seed[80],seed[1735],seed[1263],seed[1733],seed[3240],seed[3001],seed[3711],seed[741],seed[3729],seed[1550],seed[3958],seed[41],seed[348],seed[276],seed[1752],seed[2034],seed[2958],seed[996],seed[3305],seed[1162],seed[3751],seed[308],seed[1474],seed[1218],seed[920],seed[2702],seed[1755],seed[720],seed[4046],seed[3252],seed[2181],seed[2693],seed[3877],seed[2391],seed[1961],seed[1152],seed[2454],seed[1373],seed[2699],seed[1251],seed[1888],seed[1065],seed[1951],seed[659],seed[3530],seed[3113],seed[2488],seed[1751],seed[685],seed[2332],seed[3798],seed[1976],seed[2479],seed[2296],seed[1086],seed[3049],seed[2684],seed[1556],seed[597],seed[3006],seed[3464],seed[684],seed[1053],seed[3511],seed[3053],seed[1404],seed[2814],seed[3444],seed[3882],seed[542],seed[1189],seed[2623],seed[3834],seed[2727],seed[1313],seed[239],seed[3506],seed[1172],seed[3146],seed[2771],seed[1211],seed[4040],seed[3043],seed[640],seed[1322],seed[2541],seed[2245],seed[2373],seed[77],seed[1192],seed[2491],seed[2424],seed[3983],seed[2995],seed[477],seed[3483],seed[360],seed[679],seed[3914],seed[2879],seed[4041],seed[402],seed[1683],seed[2315],seed[1695],seed[2182],seed[2946],seed[3420],seed[1345],seed[1748],seed[2030],seed[3368],seed[3552],seed[2400],seed[3964],seed[2556],seed[3932],seed[2658],seed[957],seed[2665],seed[3021],seed[3928],seed[4011],seed[3823],seed[3629],seed[1057],seed[1063],seed[3459],seed[2732],seed[1741],seed[153],seed[1538],seed[1271],seed[1999],seed[2063],seed[2961],seed[1249],seed[3376],seed[3681],seed[2524],seed[2519],seed[2284]}; 
//        seed16 <= {seed[1635],seed[1248],seed[3787],seed[2981],seed[3708],seed[1658],seed[331],seed[2234],seed[3108],seed[572],seed[2986],seed[2698],seed[878],seed[2237],seed[2413],seed[375],seed[3458],seed[3375],seed[3565],seed[525],seed[778],seed[2010],seed[136],seed[3235],seed[503],seed[505],seed[2887],seed[3699],seed[1999],seed[377],seed[1526],seed[3019],seed[3343],seed[2770],seed[2160],seed[1362],seed[2650],seed[3276],seed[3230],seed[4066],seed[731],seed[3619],seed[3483],seed[1798],seed[1187],seed[1971],seed[1638],seed[3579],seed[2028],seed[1790],seed[2992],seed[1889],seed[3764],seed[1218],seed[2086],seed[2289],seed[3029],seed[3963],seed[614],seed[1384],seed[56],seed[1239],seed[1927],seed[1315],seed[1996],seed[1656],seed[3988],seed[2186],seed[1757],seed[246],seed[3612],seed[2632],seed[3778],seed[2282],seed[3297],seed[3937],seed[3053],seed[2674],seed[1848],seed[271],seed[452],seed[2714],seed[1690],seed[1486],seed[803],seed[3745],seed[5],seed[3463],seed[1314],seed[2164],seed[3595],seed[283],seed[3114],seed[2032],seed[850],seed[686],seed[3613],seed[3071],seed[120],seed[3581],seed[2097],seed[2260],seed[490],seed[985],seed[3265],seed[711],seed[3119],seed[1318],seed[3357],seed[3869],seed[1069],seed[1832],seed[2124],seed[3540],seed[4067],seed[2216],seed[581],seed[193],seed[119],seed[1223],seed[796],seed[2339],seed[1051],seed[2752],seed[499],seed[388],seed[4087],seed[311],seed[1551],seed[52],seed[1351],seed[588],seed[3913],seed[1493],seed[994],seed[573],seed[2267],seed[1340],seed[1254],seed[4077],seed[223],seed[3634],seed[4094],seed[3130],seed[3487],seed[2795],seed[3608],seed[1843],seed[3720],seed[1725],seed[1302],seed[1027],seed[1091],seed[1780],seed[3317],seed[81],seed[1162],seed[1045],seed[1079],seed[2743],seed[354],seed[1453],seed[2620],seed[1095],seed[862],seed[2584],seed[2964],seed[1370],seed[2570],seed[1772],seed[1730],seed[2358],seed[1577],seed[1781],seed[433],seed[2672],seed[3022],seed[1132],seed[4090],seed[2299],seed[960],seed[1886],seed[2680],seed[172],seed[1936],seed[555],seed[1116],seed[884],seed[2851],seed[1164],seed[1760],seed[607],seed[3982],seed[467],seed[2214],seed[4095],seed[398],seed[1582],seed[2587],seed[4064],seed[3694],seed[501],seed[2198],seed[3045],seed[3942],seed[3006],seed[2611],seed[3650],seed[1066],seed[1192],seed[387],seed[123],seed[1785],seed[86],seed[2499],seed[892],seed[2170],seed[3417],seed[1661],seed[2586],seed[2720],seed[254],seed[84],seed[1673],seed[2852],seed[3460],seed[2573],seed[3295],seed[3548],seed[836],seed[1020],seed[3628],seed[1716],seed[767],seed[3706],seed[2490],seed[2251],seed[882],seed[2244],seed[205],seed[2414],seed[3426],seed[3534],seed[1035],seed[3535],seed[1783],seed[113],seed[1859],seed[1058],seed[3283],seed[845],seed[3233],seed[2205],seed[1731],seed[2196],seed[421],seed[2412],seed[986],seed[2129],seed[2889],seed[1699],seed[1953],seed[2641],seed[45],seed[3657],seed[187],seed[4084],seed[1556],seed[3921],seed[1289],seed[1853],seed[357],seed[2759],seed[510],seed[3396],seed[683],seed[54],seed[126],seed[911],seed[821],seed[1763],seed[2336],seed[832],seed[695],seed[3618],seed[1436],seed[2746],seed[3399],seed[999],seed[1806],seed[3365],seed[3444],seed[2772],seed[905],seed[1010],seed[1256],seed[3394],seed[628],seed[195],seed[2962],seed[3476],seed[2232],seed[1237],seed[780],seed[1378],seed[2163],seed[1086],seed[913],seed[1748],seed[544],seed[828],seed[3892],seed[2043],seed[4009],seed[2295],seed[2566],seed[2017],seed[2554],seed[958],seed[644],seed[1601],seed[275],seed[3563],seed[649],seed[730],seed[2622],seed[1286],seed[2931],seed[3035],seed[3205],seed[1574],seed[3782],seed[346],seed[2471],seed[3146],seed[265],seed[760],seed[1134],seed[1932],seed[1046],seed[988],seed[540],seed[799],seed[917],seed[3829],seed[3267],seed[3600],seed[1458],seed[3739],seed[1398],seed[889],seed[668],seed[1135],seed[3187],seed[3137],seed[2204],seed[276],seed[1878],seed[1594],seed[2423],seed[2215],seed[1048],seed[613],seed[333],seed[2476],seed[3088],seed[3727],seed[923],seed[834],seed[1750],seed[531],seed[1367],seed[3939],seed[1161],seed[1459],seed[2923],seed[2785],seed[3496],seed[975],seed[3896],seed[2046],seed[1296],seed[3559],seed[787],seed[696],seed[2099],seed[1965],seed[2426],seed[2676],seed[2758],seed[497],seed[238],seed[1136],seed[3202],seed[488],seed[1720],seed[2395],seed[79],seed[2877],seed[895],seed[2867],seed[4025],seed[396],seed[1404],seed[3587],seed[2767],seed[2876],seed[1814],seed[1963],seed[3387],seed[3450],seed[3339],seed[2217],seed[3440],seed[2734],seed[1955],seed[3503],seed[473],seed[1677],seed[1073],seed[1882],seed[3799],seed[3314],seed[2303],seed[3725],seed[1924],seed[1609],seed[838],seed[2292],seed[437],seed[2451],seed[1715],seed[179],seed[2769],seed[1964],seed[738],seed[3260],seed[2799],seed[2835],seed[3515],seed[529],seed[125],seed[873],seed[247],seed[2252],seed[3875],seed[1407],seed[763],seed[3853],seed[3076],seed[2357],seed[3116],seed[1726],seed[1316],seed[2559],seed[543],seed[2280],seed[1081],seed[3555],seed[2172],seed[817],seed[3121],seed[347],seed[2970],seed[439],seed[993],seed[3794],seed[1190],seed[2737],seed[1614],seed[941],seed[3354],seed[73],seed[1209],seed[192],seed[2229],seed[3118],seed[826],seed[3907],seed[3574],seed[3656],seed[2858],seed[9],seed[164],seed[3964],seed[2812],seed[3194],seed[3030],seed[1533],seed[2624],seed[422],seed[129],seed[1445],seed[1560],seed[1349],seed[4079],seed[514],seed[4003],seed[3471],seed[368],seed[2527],seed[3768],seed[1007],seed[3277],seed[520],seed[3944],seed[1155],seed[4054],seed[606],seed[1664],seed[761],seed[229],seed[3220],seed[2513],seed[3929],seed[3226],seed[1800],seed[3959],seed[3724],seed[587],seed[1115],seed[4033],seed[1683],seed[1366],seed[3887],seed[3732],seed[1973],seed[4030],seed[3920],seed[1252],seed[719],seed[1185],seed[62],seed[4020],seed[3954],seed[807],seed[3500],seed[105],seed[1053],seed[1562],seed[944],seed[3814],seed[1128],seed[269],seed[2391],seed[2958],seed[3228],seed[815],seed[1692],seed[1172],seed[1326],seed[2219],seed[3897],seed[1666],seed[626],seed[3298],seed[1141],seed[3624],seed[2512],seed[2440],seed[2702],seed[3863],seed[1672],seed[2987],seed[1186],seed[771],seed[2464],seed[1383],seed[2274],seed[380],seed[2265],seed[2226],seed[2128],seed[3854],seed[1849],seed[3900],seed[1280],seed[3777],seed[1842],seed[2177],seed[946],seed[2056],seed[237],seed[3224],seed[1758],seed[3025],seed[487],seed[1345],seed[1625],seed[2115],seed[1472],seed[2757],seed[1344],seed[485],seed[3369],seed[177],seed[535],seed[2338],seed[3512],seed[617],seed[2378],seed[2728],seed[3360],seed[493],seed[1628],seed[3358],seed[3607],seed[457],seed[1338],seed[2488],seed[14],seed[933],seed[3598],seed[1201],seed[3684],seed[2509],seed[2319],seed[635],seed[1586],seed[3451],seed[3181],seed[3752],seed[1468],seed[3304],seed[527],seed[3240],seed[1225],seed[257],seed[1928],seed[3805],seed[1301],seed[4032],seed[1153],seed[1629],seed[2293],seed[964],seed[679],seed[255],seed[4076],seed[3553],seed[1452],seed[2318],seed[227],seed[833],seed[3385],seed[2917],seed[3832],seed[2550],seed[1372],seed[2626],seed[3671],seed[2397],seed[1170],seed[500],seed[2556],seed[1166],seed[1630],seed[848],seed[2606],seed[1513],seed[3625],seed[1102],seed[1159],seed[2246],seed[3957],seed[3253],seed[3986],seed[2079],seed[3946],seed[1126],seed[3893],seed[1967],seed[2685],seed[829],seed[1015],seed[3824],seed[441],seed[3316],seed[1188],seed[3672],seed[3315],seed[1455],seed[1534],seed[2571],seed[75],seed[181],seed[608],seed[2315],seed[1087],seed[1401],seed[3131],seed[2988],seed[2057],seed[1142],seed[2891],seed[1064],seed[2808],seed[1013],seed[3701],seed[2409],seed[2740],seed[1481],seed[218],seed[618],seed[2220],seed[3862],seed[3651],seed[1558],seed[843],seed[3482],seed[656],seed[1580],seed[290],seed[1879],seed[1307],seed[2590],seed[1568],seed[1382],seed[11],seed[4016],seed[2820],seed[224],seed[585],seed[849],seed[1516],seed[3427],seed[2106],seed[3423],seed[1129],seed[3027],seed[3132],seed[1437],seed[3830],seed[3322],seed[2258],seed[3686],seed[4024],seed[1778],seed[2594],seed[26],seed[3643],seed[3207],seed[2257],seed[855],seed[1423],seed[2608],seed[2742],seed[138],seed[330],seed[3580],seed[3851],seed[2083],seed[676],seed[2472],seed[2037],seed[1840],seed[2076],seed[3200],seed[1868],seed[3902],seed[3028],seed[447],seed[394],seed[660],seed[2657],seed[1290],seed[629],seed[2662],seed[3032],seed[1418],seed[270],seed[423],seed[942],seed[1828],seed[1341],seed[1396],seed[3812],seed[2788],seed[1575],seed[1305],seed[2779],seed[2192],seed[689],seed[579],seed[1475],seed[3818],seed[171],seed[2535],seed[3052],seed[2422],seed[2569],seed[2363],seed[2450],seed[1055],seed[2784],seed[3308],seed[2277],seed[2739],seed[3134],seed[2792],seed[1976],seed[2644],seed[3804],seed[4078],seed[3537],seed[2209],seed[3713],seed[1665],seed[3962],seed[1805],seed[2410],seed[463],seed[3871],seed[1706],seed[3721],seed[1520],seed[64],seed[3243],seed[1860],seed[1460],seed[1782],seed[2651],seed[1968],seed[1959],seed[321],seed[1917],seed[2633],seed[2848],seed[3642],seed[1031],seed[4083],seed[36],seed[996],seed[1641],seed[2945],seed[399],seed[2989],seed[3980],seed[442],seed[2883],seed[2369],seed[3860],seed[3161],seed[3345],seed[260],seed[812],seed[720],seed[819],seed[1392],seed[2591],seed[2582],seed[2560],seed[3278],seed[306],seed[2195],seed[2922],seed[3857],seed[1866],seed[918],seed[610],seed[1517],seed[2839],seed[1266],seed[4056],seed[411],seed[557],seed[1264],seed[2558],seed[1913],seed[1844],seed[3926],seed[160],seed[3490],seed[728],seed[3592],seed[2469],seed[2080],seed[2530],seed[340],seed[2806],seed[1737],seed[464],seed[3227],seed[2415],seed[1371],seed[1143],seed[222],seed[3184],seed[2328],seed[1637],seed[1273],seed[847],seed[1532],seed[402],seed[1105],seed[1140],seed[1283],seed[2087],seed[2311],seed[1705],seed[1989],seed[3763],seed[1240],seed[198],seed[2240],seed[1179],seed[870],seed[3178],seed[758],seed[3825],seed[2996],seed[3519],seed[1538],seed[2343],seed[3705],seed[3185],seed[939],seed[496],seed[672],seed[742],seed[1108],seed[1617],seed[1449],seed[153],seed[1678],seed[2640],seed[3311],seed[3372],seed[400],seed[846],seed[777],seed[2718],seed[3941],seed[1009],seed[2661],seed[2896],seed[3293],seed[2747],seed[703],seed[1138],seed[1297],seed[665],seed[1160],seed[363],seed[3556],seed[1242],seed[3631],seed[1738],seed[2437],seed[59],seed[2007],seed[1230],seed[2899],seed[3873],seed[282],seed[943],seed[3401],seed[2932],seed[1040],seed[3326],seed[1462],seed[3649],seed[978],seed[2176],seed[646],seed[2929],seed[2663],seed[1361],seed[3468],seed[391],seed[85],seed[190],seed[2143],seed[2998],seed[997],seed[3397],seed[813],seed[3215],seed[664],seed[2952],seed[3279],seed[3213],seed[3648],seed[3952],seed[3481],seed[511],seed[2646],seed[677],seed[1523],seed[185],seed[2365],seed[3973],seed[2960],seed[699],seed[2392],seed[317],seed[1615],seed[1885],seed[3232],seed[3470],seed[3066],seed[4089],seed[2436],seed[274],seed[2121],seed[2230],seed[3198],seed[3049],seed[981],seed[132],seed[2404],seed[3918],seed[2708],seed[1888],seed[4072],seed[623],seed[1946],seed[2921],seed[66],seed[1415],seed[1691],seed[1529],seed[1986],seed[453],seed[3390],seed[3932],seed[3433],seed[1576],seed[3856],seed[1454],seed[3239],seed[252],seed[1395],seed[1060],seed[2555],seed[3912],seed[2323],seed[1792],seed[4007],seed[3802],seed[3204],seed[995],seed[2713],seed[1113],seed[2879],seed[3211],seed[359],seed[448],seed[1605],seed[823],seed[897],seed[2574],seed[3036],seed[1700],seed[2557],seed[1708],seed[197],seed[3806],seed[558],seed[3521],seed[955],seed[3465],seed[3415],seed[4039],seed[797],seed[2025],seed[147],seed[3009],seed[3575],seed[934],seed[3868],seed[512],seed[1773],seed[1090],seed[4069],seed[2459],seed[2045],seed[2704],seed[559],seed[1646],seed[2701],seed[3425],seed[1648],seed[2592],seed[3325],seed[725],seed[209],seed[1569],seed[292],seed[1542],seed[2071],seed[3095],seed[3928],seed[2690],seed[2968],seed[3165],seed[1123],seed[1310],seed[3400],seed[3557],seed[3828],seed[974],seed[443],seed[3186],seed[2144],seed[1775],seed[2859],seed[1680],seed[2589],seed[3916],seed[1825],seed[1890],seed[1306],seed[3743],seed[984],seed[586],seed[3518],seed[876],seed[2073],seed[1385],seed[3176],seed[2107],seed[3827],seed[1815],seed[2145],seed[41],seed[1549],seed[1626],seed[2496],seed[1983],seed[4037],seed[3590],seed[2110],seed[582],seed[1940],seed[2673],seed[3632],seed[3622],seed[1279],seed[3287],seed[2473],seed[1444],seed[2810],seed[3193],seed[1198],seed[1098],seed[3975],seed[701],seed[2201],seed[602],seed[2432],seed[3418],seed[2354],seed[1016],seed[2683],seed[2818],seed[2278],seed[3138],seed[1537],seed[3381],seed[1883],seed[1813],seed[899],seed[3785],seed[998],seed[407],seed[2925],seed[1528],seed[3229],seed[2732],seed[80],seed[810],seed[2462],seed[1085],seed[861],seed[3620],seed[783],seed[1573],seed[1291],seed[2390],seed[630],seed[970],seed[3175],seed[3145],seed[2006],seed[888],seed[2933],seed[1590],seed[1078],seed[3439],seed[2327],seed[1911],seed[3583],seed[1751],seed[1490],seed[1662],seed[1521],seed[3728],seed[72],seed[502],seed[343],seed[2030],seed[1104],seed[47],seed[2763],seed[1717],seed[1689],seed[2340],seed[2572],seed[2285],seed[1793],seed[1922],seed[1564],seed[1446],seed[2712],seed[908],seed[3577],seed[2607],seed[118],seed[371],seed[281],seed[2817],seed[2865],seed[416],seed[2691],seed[1895],seed[3221],seed[2502],seed[3610],seed[1548],seed[3864],seed[325],seed[2184],seed[616],seed[1695],seed[710],seed[3442],seed[2537],seed[1281],seed[4010],seed[2202],seed[3816],seed[1795],seed[2719],seed[2168],seed[764],seed[2609],seed[3726],seed[1624],seed[1912],seed[355],seed[980],seed[251],seed[1410],seed[2872],seed[2565],seed[662],seed[621],seed[1246],seed[3323],seed[1313],seed[3978],seed[1257],seed[3850],seed[3955],seed[174],seed[294],seed[605],seed[3740],seed[1364],seed[3395],seed[3309],seed[1175],seed[2910],seed[3508],seed[3710],seed[3709],seed[3301],seed[1325],seed[3539],seed[2302],seed[4],seed[2181],seed[3270],seed[2048],seed[576],seed[4045],seed[53],seed[207],seed[3582],seed[2297],seed[563],seed[781],seed[3344],seed[979],seed[2016],seed[3231],seed[87],seed[948],seed[2012],seed[320],seed[2829],seed[1740],seed[1707],seed[4029],seed[1334],seed[2652],seed[3303],seed[83],seed[2372],seed[1687],seed[1839],seed[1150],seed[454],seed[1319],seed[3330],seed[762],seed[3754],seed[465],seed[2900],seed[2744],seed[3822],seed[2194],seed[184],seed[2489],seed[3685],seed[2705],seed[3536],seed[2875],seed[2287],seed[3691],seed[3605],seed[1328],seed[1583],seed[1921],seed[1089],seed[3441],seed[3434],seed[250],seed[1704],seed[1514],seed[2250],seed[1933],seed[740],seed[3562],seed[1835],seed[0],seed[3288],seed[3089],seed[1269],seed[2005],seed[176],seed[2729],seed[298],seed[713],seed[3674],seed[792],seed[3333],seed[322],seed[3588],seed[3275],seed[2162],seed[3180],seed[3000],seed[2627],seed[1919],seed[611],seed[2174],seed[3696],seed[1251],seed[4012],seed[1623],seed[2508],seed[3846],seed[3569],seed[2070],seed[2088],seed[1434],seed[2157],seed[1891],seed[300],seed[3561],seed[519],seed[428],seed[2974],seed[2761],seed[3596],seed[1465],seed[2724],seed[3750],seed[2826],seed[2183],seed[1747],seed[2361],seed[3],seed[384],seed[358],seed[432],seed[1125],seed[3210],seed[1610],seed[1375],seed[2382],seed[1612],seed[3452],seed[2679],seed[3190],seed[1387],seed[3773],seed[580],seed[3578],seed[1097],seed[3981],seed[2881],seed[312],seed[2843],seed[914],seed[2134],seed[1299],seed[2261],seed[1650],seed[1771],seed[3905],seed[3154],seed[989],seed[2091],seed[734],seed[3015],seed[2044],seed[702],seed[1915],seed[2453],seed[3256],seed[2228],seed[173],seed[6],seed[1600],seed[2693],seed[1808],seed[1212],seed[291],seed[4026],seed[178],seed[3718],seed[750],seed[2773],seed[1850],seed[309],seed[3044],seed[3621],seed[134],seed[263],seed[3192],seed[121],seed[97],seed[264],seed[1694],seed[3408],seed[2098],seed[3584],seed[3055],seed[2478],seed[2920],seed[2643],seed[33],seed[2275],seed[1106],seed[2135],seed[2367],seed[3173],seed[2903],seed[3516],seed[612],seed[2018],seed[124],seed[3447],seed[338],seed[2101],seed[652],seed[1033],seed[2094],seed[1036],seed[1743],seed[1137],seed[3693],seed[2222],seed[1011],seed[3938],seed[1670],seed[1380],seed[3550],seed[3477],seed[1987],seed[3765],seed[2360],seed[2428],seed[2002],seed[953],seed[3082],seed[2616],seed[3646],seed[1505],seed[2790],seed[3532],seed[2371],seed[1916],seed[3286],seed[2211],seed[2778],seed[3876],seed[418],seed[2435],seed[2465],seed[3993],seed[739],seed[1755],seed[3925],seed[2575],seed[2114],seed[504],seed[1711],seed[756],seed[1768],seed[2189],seed[3453],seed[25],seed[2534],seed[2515],seed[1535],seed[2653],seed[1145],seed[3046],seed[2975],seed[1061],seed[3112],seed[3072],seed[726],seed[2544],seed[3527],seed[2716],seed[1657],seed[765],seed[1466],seed[3927],seed[1093],seed[1567],seed[383],seed[2993],seed[1205],seed[2380],seed[3206],seed[3282],seed[2449],seed[492],seed[2431],seed[356],seed[1496],seed[3554],seed[372],seed[3617],seed[2288],seed[2433],seed[1381],seed[189],seed[522],seed[3247],seed[3826],seed[2581],seed[2617],seed[1647],seed[2904],seed[150],seed[151],seed[1679],seed[1447],seed[1732],seed[1259],seed[3086],seed[494],seed[3012],seed[539],seed[1881],seed[3241],seed[2748],seed[3337],seed[794],seed[3681],seed[716],seed[655],seed[2760],seed[4014],seed[2480],seed[589],seed[3122],seed[3169],seed[1030],seed[1443],seed[2294],seed[3890],seed[2182],seed[3984],seed[650],seed[3786],seed[3329],seed[2798],seed[2520],seed[1676],seed[2350],seed[2103],seed[2347],seed[3371],seed[4086],seed[2601],seed[1063],seed[1482],seed[2501],seed[2169],seed[455],seed[3769],seed[2655],seed[231],seed[2753],seed[3968],seed[484],seed[951],seed[2786],seed[546],seed[3074],seed[4046],seed[2159],seed[459],seed[566],seed[2377],seed[3430],seed[3711],seed[2486],seed[395],seed[155],seed[3811],seed[2063],seed[1993],seed[3429],seed[68],seed[1037],seed[1285],seed[3910],seed[1471],seed[2963],seed[140],seed[145],seed[3081],seed[1620],seed[2782],seed[3380],seed[2949],seed[789],seed[2504],seed[406],seed[95],seed[3140],seed[775],seed[288],seed[1148],seed[1803],seed[3623],seed[568],seed[1884],seed[2972],seed[2061],seed[2855],seed[3498],seed[1207],seed[2514],seed[1429],seed[2816],seed[2831],seed[1876],seed[2495],seed[2364],seed[2938],seed[74],seed[601],seed[1421],seed[3393],seed[596],seed[3179],seed[1831],seed[4013],seed[1962],seed[3652],seed[3378],seed[1602],seed[1473],seed[1502],seed[688],seed[1425],seed[1109],seed[2600],seed[1960],seed[749],seed[2588],seed[35],seed[3790],seed[722],seed[3334],seed[3741],seed[2510],seed[3940],seed[3064],seed[2888],seed[1497],seed[506],seed[1177],seed[2916],seed[272],seed[2402],seed[3174],seed[909],seed[1863],seed[1117],seed[89],seed[3057],seed[1920],seed[3070],seed[1197],seed[1952],seed[1184],seed[285],seed[3915],seed[1599],seed[1287],seed[2541],seed[3586],seed[793],seed[71],seed[382],seed[2847],seed[1833],seed[1943],seed[3712],seed[2188],seed[3560],seed[201],seed[3300],seed[1193],seed[3061],seed[746],seed[410],seed[415],seed[2411],seed[1320],seed[1561],seed[2796],seed[3966],seed[1898],seed[4038],seed[133],seed[2154],seed[3110],seed[2055],seed[3100],seed[91],seed[213],seed[2854],seed[65],seed[3788],seed[3488],seed[1120],seed[1413],seed[2730],seed[1552],seed[1167],seed[3517],seed[1288],seed[361],seed[3636],seed[654],seed[390],seed[3819],seed[1622],seed[2109],seed[1801],seed[3217],seed[3789],seed[1820],seed[2850],seed[1660],seed[1713],seed[16],seed[3435],seed[600],seed[3336],seed[348],seed[2000],seed[3965],seed[2457],seed[217],seed[2379],seed[1356],seed[1448],seed[2393],seed[3250],seed[1937],seed[1216],seed[2036],seed[1788],seed[426],seed[1270],seed[339],seed[2108],seed[2003],seed[2642],seed[4088],seed[4055],seed[3058],seed[2243],seed[3328],seed[2648],seed[2985],seed[1871],seed[2546],seed[3269],seed[3771],seed[2033],seed[3775],seed[3678],seed[865],seed[3109],seed[2112],seed[3416],seed[3813],seed[1598],seed[2286],seed[2042],seed[2678],seed[3382],seed[3263],seed[867],seed[2041],seed[1337],seed[161],seed[1753],seed[130],seed[2551],seed[3364],seed[2474],seed[3424],seed[2466],seed[1817],seed[2381],seed[1094],seed[3376],seed[3107],seed[3411],seed[801],seed[592],seed[1227],seed[2756],seed[881],seed[2139],seed[3502],seed[144],seed[2349],seed[1154],seed[2305],seed[859],seed[3274],seed[1034],seed[3048],seed[477],seed[3523],seed[3341],seed[2062],seed[634],seed[1202],seed[2579],seed[550],seed[3351],seed[3606],seed[732],seed[1746],seed[214],seed[1477],seed[3974],seed[4031],seed[2346],seed[864],seed[3128],seed[2687],seed[3983],seed[2629],seed[1234],seed[1304],seed[643],seed[2482],seed[2997],seed[860],seed[903],seed[77],seed[4047],seed[2445],seed[374],seed[169],seed[2442],seed[2052],seed[3105],seed[3037],seed[3919],seed[1492],seed[837],seed[1530],seed[1544],seed[3111],seed[3914],seed[1054],seed[3356],seed[1335],seed[2863],seed[3246],seed[3703],seed[2539],seed[2040],seed[3770],seed[1830],seed[3970],seed[2545],seed[305],seed[2038],seed[2383],seed[1565],seed[715],seed[329],seed[1988],seed[163],seed[2707],seed[1938],seed[3238],seed[2291],seed[32],seed[3747],seed[1906],seed[27],seed[2241],seed[2264],seed[670],seed[1893],seed[3492],seed[168],seed[2185],seed[1480],seed[3059],seed[3366],seed[232],seed[1494],seed[2549],seed[2621],seed[1461],seed[239],seed[751],seed[532],seed[3189],seed[690],seed[1697],seed[717],seed[1518],seed[2517],seed[4063],seed[3735],seed[827],seed[904],seed[3342],seed[444],seed[2425],seed[3249],seed[3697],seed[3865],seed[3318],seed[3626],seed[2930],seed[1762],seed[1639],seed[1284],seed[627],seed[2822],seed[3023],seed[3729],seed[3063],seed[647],seed[542],seed[2647],seed[1408],seed[2446],seed[2950],seed[2585],seed[324],seed[3151],seed[795],seed[2577],seed[2253],seed[491],seed[2388],seed[3248],seed[3738],seed[2825],seed[929],seed[4035],seed[2834],seed[167],seed[1634],seed[1438],seed[2254],seed[2543],seed[1004],seed[2861],seed[127],seed[3704],seed[645],seed[381],seed[3234],seed[2866],seed[2179],seed[3486],seed[2353],seed[3414],seed[1228],seed[2856],seed[1232],seed[3080],seed[2193],seed[641],seed[370],seed[3043],seed[3670],seed[3664],seed[4091],seed[661],seed[2604],seed[874],seed[1826],seed[822],seed[1277],seed[15],seed[1804],seed[1642],seed[1651],seed[157],seed[435],seed[3493],seed[1539],seed[2213],seed[3142],seed[3667],seed[620],seed[2065],seed[755],seed[3011],seed[2631],seed[2765],seed[533],seed[2366],seed[293],seed[3855],seed[1742],seed[2078],seed[1017],seed[3753],seed[1439],seed[2635],seed[1770],seed[2406],seed[413],seed[2939],seed[3969],seed[3067],seed[456],seed[3541],seed[1139],seed[3075],seed[685],seed[3715],seed[1794],seed[536],seed[3096],seed[2552],seed[785],seed[3117],seed[1261],seed[2148],seed[2419],seed[1718],seed[3679],seed[2967],seed[940],seed[2871],seed[651],seed[2845],seed[2484],seed[1873],seed[1221],seed[2180],seed[3604],seed[830],seed[1243],seed[3707],seed[1767],seed[3630],seed[2598],seed[1531],seed[2105],seed[475],seed[2892],seed[707],seed[2069],seed[462],seed[2966],seed[2731],seed[952],seed[1945],seed[3756],seed[2942],seed[1616],seed[2941],seed[3934],seed[2004],seed[3682],seed[3861],seed[741],seed[1667],seed[13],seed[2092],seed[7],seed[2522],seed[1379],seed[624],seed[341],seed[3195],seed[335],seed[2421],seed[2191],seed[262],seed[244],seed[3525],seed[1925],seed[959],seed[3445],seed[342],seed[2399],seed[1816],seed[2233],seed[3284],seed[3392],seed[615],seed[2727],seed[3047],seed[420],seed[637],seed[1595],seed[2959],seed[3412],seed[1350],seed[3148],seed[1961],seed[2138],seed[2533],seed[1038],seed[947],seed[1183],seed[267],seed[2983],seed[3638],seed[3666],seed[1607],seed[191],seed[3877],seed[1572],seed[2123],seed[2256],seed[3759],seed[286],seed[2531],seed[1321],seed[3324],seed[3923],seed[1099],seed[3079],seed[3144],seed[3362],seed[2971],seed[438],seed[3979],seed[3398],seed[3662],seed[852],seed[2368],seed[737],seed[1969],seed[364],seed[1649],seed[2085],seed[574],seed[3888],seed[991],seed[820],seed[1426],seed[1511],seed[636],seed[774],seed[2334],seed[3355],seed[3884],seed[3348],seed[591],seed[1908],seed[2218],seed[3641],seed[1579],seed[3428],seed[2807],seed[352],seed[2681],seed[928],seed[2460],seed[3616],seed[1047],seed[3335],seed[3281],seed[2776],seed[3251],seed[1698],seed[3242],seed[48],seed[334],seed[3403],seed[2401],seed[3208],seed[609],seed[102],seed[2141],seed[389],seed[4036],seed[2862],seed[3083],seed[1627],seed[2783],seed[1399],seed[1174],seed[2583],seed[3528],seed[3924],seed[3901],seed[2269],seed[1684],seed[1734],seed[3084],seed[3489],seed[2630],seed[2122],seed[3796],seed[1841],seed[2936],seed[3338],seed[307],seed[3219],seed[3717],seed[759],seed[863],seed[1491],seed[109],seed[773],seed[2394],seed[2529],seed[2605],seed[1057],seed[570],seed[3160],seed[4041],seed[3222],seed[2692],seed[1929],seed[3167],seed[2781],seed[2578],seed[78],seed[2898],seed[2658],seed[412],seed[2456],seed[3762],seed[2821],seed[2519],seed[1702],seed[3820],seed[2645],seed[3257],seed[3730],seed[373],seed[3158],seed[3254],seed[508],seed[898],seed[3102],seed[297],seed[3010],seed[3272],seed[2787],seed[2084],seed[1709],seed[3629],seed[3368],seed[2116],seed[1092],seed[104],seed[3858],seed[631],seed[1268],seed[3766],seed[2722],seed[806],seed[1008],seed[2072],seed[57],seed[3018],seed[2666],seed[976],seed[1581],seed[2498],seed[1724],seed[3698],seed[1478],seed[598],seed[1838],seed[1176],seed[2823],seed[3669],seed[3472],seed[2173],seed[3776],seed[2344],seed[2384],seed[1896],seed[2800],seed[2766],seed[107],seed[2842],seed[2444],seed[3835],seed[927],seed[3410],seed[234],seed[2161],seed[1352],seed[3683],seed[1653],seed[745],seed[2326],seed[1430],seed[3021],seed[551],seed[3882],seed[3842],seed[3040],seed[887],seed[2126],seed[3880],seed[2373],seed[957],seed[2166],seed[1631],seed[4050],seed[809],seed[1809],seed[2492],seed[3947],seed[1376],seed[2567],seed[2470],seed[3594],seed[2111],seed[1741],seed[1411],seed[3172],seed[642],seed[3259],seed[2307],seed[1854],seed[1433],seed[3599],seed[1072],seed[1118],seed[367],seed[204],seed[1181],seed[790],seed[961],seed[1857],seed[3639],seed[965],seed[2723],seed[1278],seed[916],seed[2158],seed[886],seed[680],seed[240],seed[3404],seed[727],seed[3719],seed[2049],seed[2019],seed[1640],seed[2526],seed[779],seed[3961],seed[110],seed[4015],seed[196],seed[2247],seed[1686],seed[901],seed[4059],seed[2420],seed[2654],seed[301],seed[3383],seed[1956],seed[1173],seed[2483],seed[1761],seed[3113],seed[2832],seed[1931],seed[135],seed[2726],seed[203],seed[3386],seed[405],seed[296],seed[2775],seed[202],seed[1000],seed[128],seed[816],seed[1019],seed[2156],seed[1942],seed[414],seed[2479],seed[1180],seed[1597],seed[2675],seed[597],seed[1984],seed[2901],seed[474],seed[1133],seed[2638],seed[1059],seed[3654],seed[3520],seed[2375],seed[982],seed[137],seed[648],seed[3972],seed[2133],seed[1103],seed[2427],seed[149],seed[480],seed[3702],seed[2564],seed[2880],seed[2669],seed[851],seed[1618],seed[885],seed[386],seed[1570],seed[3748],seed[575],seed[1654],seed[1],seed[76],seed[360],seed[1902],seed[983],seed[4040],seed[3252],seed[378],seed[2059],seed[1926],seed[3737],seed[883],seed[3791],seed[1671],seed[1112],seed[3746],seed[1463],seed[1789],seed[2870],seed[1327],seed[3157],seed[2245],seed[4071],seed[2095],seed[1990],seed[924],seed[2697],seed[736],seed[55],seed[2505],seed[2058],seed[2794],seed[4018],seed[38],seed[673],seed[1200],seed[3546],seed[962],seed[34],seed[1258],seed[3558],seed[561],seed[3547],seed[3817],seed[2325],seed[2497],seed[4043],seed[450],seed[1519],seed[3191],seed[2200],seed[1723],seed[4053],seed[3031],seed[2322],seed[3307],seed[289],seed[1483],seed[2677],seed[3377],seed[43],seed[1076],seed[1196],seed[3120],seed[2239],seed[1331],seed[920],seed[3094],seed[2494],seed[593],seed[2503],seed[3742],seed[249],seed[931],seed[3576],seed[2793],seed[17],seed[1571],seed[3511],seed[3182],seed[1068],seed[2352],seed[2153],seed[2175],seed[3352],seed[1359],seed[2370],seed[4068],seed[4073],seed[1217],seed[1414],seed[2255],seed[2400],seed[2836],seed[709],seed[2348],seed[1507],seed[2356],seed[1923],seed[98],seed[1424],seed[2755],seed[1712],seed[1824],seed[3268],seed[1336],seed[3155],seed[4042],seed[3522],seed[4070],seed[2809],seed[528],seed[287],seed[2523],seed[930],seed[268],seed[3544],seed[800],seed[182],seed[1901],seed[2894],seed[2837],seed[3843],seed[3834],seed[1547],seed[2500],seed[1213],seed[2281],seed[2750],seed[1124],seed[3197],seed[2090],seed[1071],seed[228],seed[3953],seed[714],seed[2946],seed[3609],seed[3209],seed[788],seed[1950],seed[708],seed[2634],seed[482],seed[1157],seed[2104],seed[2853],seed[2660],seed[1353],seed[1215],seed[3319],seed[2051],seed[3614],seed[1644],seed[967],seed[233],seed[1122],seed[1752],seed[108],seed[1948],seed[3676],seed[1796],seed[3585],seed[3551],seed[3042],seed[3513],seed[3722],seed[362],seed[2548],seed[1722],seed[1769],seed[2403],seed[3466],seed[401],seed[115],seed[1158],seed[3549],seed[1119],seed[638],seed[22],seed[1163],seed[3886],seed[154],seed[1342],seed[1836],seed[1080],seed[3236],seed[1373],seed[3680],seed[3781],seed[1765],seed[2113],seed[2602],seed[2331],seed[3419],seed[3744],seed[4017],seed[1088],seed[1100],seed[67],seed[3420],seed[2542],seed[910],seed[2387],seed[2074],seed[2994],seed[1470],seed[2840],seed[1823],seed[3695],seed[3971],seed[1500],seed[2487],seed[1348],seed[1169],seed[857],seed[3005],seed[1555],seed[3087],seed[142],seed[1479],seed[3529],seed[3506],seed[1435],seed[1220],seed[906],seed[4057],seed[345],seed[4052],seed[2454],seed[3056],seed[554],seed[769],seed[782],seed[2937],seed[3815],seed[3153],seed[3407],seed[3289],seed[972],seed[3150],seed[3542],seed[2385],seed[3573],seed[2026],seed[2689],seed[3361],seed[1365],seed[3690],seed[772],seed[2736],seed[1970],seed[2979],seed[1357],seed[3644],seed[69],seed[4019],seed[2868],seed[1032],seed[577],seed[2203],seed[3658],seed[3568],seed[2389],seed[798],seed[417],seed[1333],seed[2068],seed[349],seed[1210],seed[489],seed[541],seed[2506],seed[971],seed[2408],seed[3602],seed[3524],seed[3196],seed[4049],seed[1875],seed[1253],seed[2667],seed[253],seed[1633],seed[302],seed[658],seed[681],seed[2308],seed[1764],seed[2637],seed[2351],seed[4060],seed[1377],seed[2027],seed[1298],seed[3688],seed[1903],seed[877],seed[2918],seed[3883],seed[2668],seed[436],seed[1587],seed[2982],seed[8],seed[2686],seed[3104],seed[2991],seed[2272],seed[3183],seed[2011],seed[365],seed[2999],seed[2948],seed[3572],seed[2165],seed[3533],seed[101],seed[1675],seed[1818],seed[814],seed[2321],seed[2022],seed[1219],seed[1543],seed[1236],seed[2398],seed[691],seed[1250],seed[839],seed[2664],seed[328],seed[1827],seed[313],seed[2429],seed[476],seed[1206],seed[2066],seed[230],seed[2117],seed[2857],seed[2849],seed[308],seed[534],seed[3784],seed[3432],seed[3212],seed[2493],seed[2467],seed[516],seed[3731],seed[578],seed[4021],seed[704],seed[460],seed[4034],seed[2738],seed[3258],seed[486],seed[752],seed[4082],seed[1862],seed[3456],seed[3168],seed[2768],seed[729],seed[2020],seed[3162],seed[3749],seed[2990],seed[1872],seed[1865],seed[376],seed[3384],seed[1503],seed[51],seed[2050],seed[1235],seed[425],seed[2485],seed[1386],seed[3845],seed[723],seed[1419],seed[804],seed[925],seed[1292],seed[2908],seed[3106],seed[256],seed[3564],seed[3917],seed[3092],seed[1525],seed[3994],seed[1312],seed[1402],seed[1802],seed[1489],seed[1696],seed[791],seed[3484],seed[199],seed[2995],seed[523],seed[3203],seed[2961],seed[220],seed[369],seed[3844],seed[2603],seed[165],seed[3216],seed[1759],seed[2093],seed[968],seed[215],seed[2481],seed[3531],seed[1632],seed[2984],seed[869],seed[2943],seed[3872],seed[2301],seed[12],seed[3767],seed[1958],seed[2670],seed[2771],seed[3346],seed[3640],seed[440],seed[3504],seed[186],seed[973],seed[2082],seed[3507],seed[1147],seed[1588],seed[2430],seed[935],seed[1189],seed[571],seed[1710],seed[3370],seed[743],seed[3809],seed[524],seed[397],seed[2407],seed[408],seed[1749],seed[2595],seed[595],seed[2314],seed[3772],seed[4093],seed[1405],seed[1897],seed[4006],seed[2568],seed[1829],seed[3894],seed[2919],seed[3285],seed[1432],seed[818],seed[2907],seed[404],seed[2711],seed[3026],seed[1861],seed[2310],seed[279],seed[3436],seed[1231],seed[211],seed[950],seed[1168],seed[332],seed[3340],seed[3388],seed[3171],seed[875],seed[1001],seed[3881],seed[1957],seed[1655],seed[42],seed[1420],seed[3007],seed[954],seed[49],seed[1596],seed[1777],seed[2873],seed[1309],seed[1146],seed[1262],seed[2780],seed[1499],seed[2897],seed[3093],seed[1563],seed[692],seed[3552],seed[2789],seed[2284],seed[166],seed[932],seed[2001],seed[2441],seed[424],seed[1247],seed[507],seed[1527],seed[1317],seed[1845],seed[3402],seed[2813],seed[2249],seed[2235],seed[3976],seed[3645],seed[1797],seed[640],seed[2935],seed[2725],seed[871],seed[3647],seed[471],seed[2553],seed[188],seed[949],seed[1974],seed[1042],seed[1211],seed[1476],seed[2562],seed[1006],seed[3099],seed[2],seed[1980],seed[1014],seed[842],seed[858],seed[560],seed[92],seed[2024],seed[2197],seed[1807],seed[2268],seed[1276],seed[1992],seed[3795],seed[556],seed[1892],seed[3462],seed[1339],seed[219],seed[2424],seed[2064],seed[114],seed[2610],seed[2227],seed[2954],seed[900],seed[1786],seed[1869],seed[2376],seed[2521],seed[19],seed[1245],seed[1224],seed[824],seed[39],seed[1997],seed[226],seed[1811],seed[1203],seed[2944],seed[1506],seed[1918],seed[2132],seed[1501],seed[2374],seed[152],seed[678],seed[3841],seed[3780],seed[3024],seed[1721],seed[1659],seed[241],seed[1776],seed[3627],seed[584],seed[2947],seed[3147],seed[3904],seed[3838],seed[1431],seed[1368],seed[1238],seed[61],seed[2869],seed[784],seed[553],seed[1899],seed[2448],seed[2015],seed[2060],seed[1084],seed[2054],seed[1604],seed[2455],seed[2309],seed[1681],seed[2150],seed[3989],seed[3320],seed[748],seed[1719],seed[1589],seed[992],seed[2953],seed[526],seed[3363],seed[3473],seed[3797],seed[1606],seed[2341],seed[4023],seed[3266],seed[3464],seed[3001],seed[3016],seed[667],seed[3313],seed[481],seed[633],seed[461],seed[4085],seed[2814],seed[1682],seed[20],seed[1272],seed[4092],seed[3996],seed[1474],seed[3421],seed[682],seed[1303],seed[3839],seed[3069],seed[537],seed[3479],seed[3133],seed[1096],seed[1263],seed[3136],seed[786],seed[3908],seed[549],seed[2864],seed[945],seed[768],seed[1566],seed[4011],seed[1856],seed[2684],seed[2119],seed[3262],seed[3933],seed[88],seed[893],seed[3758],seed[2618],seed[3332],seed[3103],seed[3950],seed[3405],seed[2271],seed[603],seed[3469],seed[2639],seed[1541],seed[2625],seed[344],seed[208],seed[3115],seed[3505],seed[2075],seed[1852],seed[379],seed[3859],seed[1578],seed[705],seed[1442],seed[2223],seed[304],seed[990],seed[1951],seed[1182],seed[2884],seed[3803],seed[143],seed[2665],seed[2804],seed[2547],seed[1979],seed[1025],seed[295],seed[2940],seed[840],seed[24],seed[1417],seed[1985],seed[3051],seed[141],seed[4008],seed[1195],seed[46],seed[1311],seed[1024],seed[1322],seed[969],seed[29],seed[2089],seed[2576],seed[2386],seed[698],seed[299],seed[754],seed[835],seed[1733],seed[112],seed[2957],seed[111],seed[323],seed[1271],seed[3261],seed[3497],seed[2342],seed[3800],seed[1495],seed[3004],seed[1075],seed[70],seed[1082],seed[117],seed[1409],seed[674],seed[3003],seed[2764],seed[2525],seed[2805],seed[2735],seed[1260],seed[3097],seed[663],seed[2199],seed[2034],seed[3459],seed[1593],seed[2882],seed[451],seed[4028],seed[802],seed[2355],seed[3457],seed[479],seed[3170],seed[706],seed[1049],seed[562],seed[757],seed[811],seed[3264],seed[1374],seed[2890],seed[1947],seed[2047],seed[3467],seed[392],seed[3761],seed[1074],seed[583],seed[1652],seed[1619],seed[2077],seed[2927],seed[3139],seed[445],seed[3977],seed[2709],seed[2803],seed[653],seed[1779],seed[2273],seed[1121],seed[175],seed[3922],seed[1510],seed[3164],seed[3736],seed[3478],seed[4065],seed[3199],seed[2615],seed[3751],seed[243],seed[4061],seed[3936],seed[1241],seed[2283],seed[619],seed[2878],seed[58],seed[1498],seed[4062],seed[1226],seed[776],seed[3878],seed[963],seed[183],seed[2096],seed[3601],seed[3327],seed[1403],seed[419],seed[733],seed[3454],seed[2827],seed[1022],seed[1880],seed[4048],seed[3991],seed[1799],seed[2841],seed[2599],seed[3987],seed[1440],seed[2695],seed[1343],seed[2536],seed[2538],seed[3906],seed[3903],seed[599],seed[2147],seed[2928],seed[3237],seed[518],seed[2008],seed[3124],seed[1701],seed[2167],seed[3949],seed[2682],seed[4058],seed[3889],seed[2035],seed[1393],seed[1728],seed[3810],seed[697],seed[3792],seed[805],seed[880],seed[2516],seed[545],seed[3389],seed[3570],seed[1978],seed[744],seed[1065],seed[1003],seed[2345],seed[1416],seed[3041],seed[659],seed[3033],seed[1021],seed[1870],seed[3480],seed[724],seed[521],seed[2874],seed[31],seed[1111],seed[564],seed[890],seed[825],seed[1944],seed[2777],seed[2741],seed[987],seed[657],seed[1427],seed[261],seed[639],seed[3495],seed[483],seed[3545],seed[116],seed[3774],seed[103],seed[3567],seed[2102],seed[1663],seed[3166],seed[3485],seed[3135],seed[3958],seed[3060],seed[2699],seed[2236],seed[2659],seed[1165],seed[148],seed[747],seed[434],seed[326],seed[2081],seed[3367],seed[3635],seed[1855],seed[1052],seed[856],seed[2337],seed[1522],seed[2619],seed[2146],seed[2561],seed[1557],seed[2023],seed[3716],seed[3945],seed[868],seed[2131],seed[1002],seed[3127],seed[1394],seed[2021],seed[3014],seed[1509],seed[3571],seed[2951],seed[2416],seed[2100],seed[2518],seed[2330],seed[2266],seed[896],seed[3948],seed[4027],seed[469],seed[1274],seed[3951],seed[1736],seed[2934],seed[277],seed[2955],seed[1819],seed[3895],seed[3373],seed[3494],seed[2009],seed[3689],seed[1467],seed[2895],seed[2248],seed[28],seed[1591],seed[1044],seed[210],seed[200],seed[1130],seed[3931],seed[1621],seed[2924],seed[1766],seed[509],seed[318],seed[1611],seed[4000],seed[1178],seed[3002],seed[3823],seed[3008],seed[3091],seed[1998],seed[1584],seed[1585],seed[2405],seed[1464],seed[632],seed[3870],seed[3757],seed[517],seed[2532],seed[1914],seed[2434],seed[1293],seed[1360],seed[1005],seed[478],seed[3760],seed[350],seed[1553],seed[1887],seed[449],seed[1194],seed[1669],seed[1067],seed[1056],seed[3413],seed[2906],seed[2811],seed[3152],seed[1039],seed[2612],seed[273],seed[2014],seed[2893],seed[922],seed[894],seed[1295],seed[3201],seed[44],seed[3597],seed[2721],seed[530],seed[2224],seed[446],seed[1127],seed[590],seed[1347],seed[316],seed[1204],seed[3530],seed[3998],seed[2140],seed[1208],seed[1592],seed[3177],seed[1949],seed[3491],seed[3296],seed[2238],seed[3218],seed[1847],seed[3848],seed[3294],seed[3409],seed[3461],seed[2976],seed[3188],seed[1688],seed[2524],seed[1012],seed[2316],seed[212],seed[938],seed[3291],seed[162],seed[3474],seed[1905],seed[3930],seed[1693],seed[122],seed[2860],seed[18],seed[1674],seed[3431],seed[353],seed[2329],seed[1485],seed[1603],seed[82],seed[1329],seed[3700],seed[1991],seed[1191],seed[1062],seed[2458],seed[2130],seed[2335],seed[3891],seed[21],seed[1546],seed[1536],seed[3347],seed[96],seed[3125],seed[2844],seed[2306],seed[2791],seed[3141],seed[687],seed[1400],seed[3455],seed[4005],seed[4001],seed[3603],seed[1441],seed[1954],seed[1275],seed[3956],seed[1645],seed[3017],seed[3290],seed[1144],seed[2902],seed[3312],seed[1977],seed[3223],seed[225],seed[2802],seed[3911],seed[2700],seed[569],seed[3306],seed[2029],seed[3849],seed[1877],seed[4044],seed[242],seed[3543],seed[3615],seed[498],seed[3526],seed[1043],seed[3050],seed[3867],seed[2913],seed[468],seed[1214],seed[2317],seed[2715],seed[936],seed[2152],seed[259],seed[3509],seed[2563],seed[3733],seed[1981],seed[1995],seed[3292],seed[3899],seed[3078],seed[2438],seed[3663],seed[1791],seed[1834],seed[1456],seed[303],seed[2067],seed[1907],seed[2819],seed[327],seed[1735],seed[3475],seed[1643],seed[2118],seed[2828],seed[3273],seed[3831],seed[2540],seed[146],seed[712],seed[1488],seed[1041],seed[669],seed[236],seed[248],seed[4004],seed[472],seed[3065],seed[385],seed[3591],seed[3159],seed[63],seed[966],seed[10],seed[3422],seed[2149],seed[3734],seed[3349],seed[3038],seed[2231],seed[1324],seed[2210],seed[2362],seed[1982],seed[2751],seed[565],seed[1487],seed[666],seed[2797],seed[2905],seed[3156],seed[2333],seed[1323],seed[180],seed[891],seed[1972],seed[3149],seed[100],seed[770],seed[2262],seed[1894],seed[2477],seed[515],seed[3310],seed[1837],seed[1821],seed[1756],seed[2511],seed[3837],seed[1774],seed[1874],seed[3999],seed[1504],seed[1934],seed[1222],seed[3244],seed[1812],seed[4075],seed[3245],seed[1114],seed[1975],seed[2270],seed[3446],seed[2694],seed[1966],seed[194],seed[1822],seed[2909],seed[158],seed[23],seed[2463],seed[3985],seed[3593],seed[1484],seed[221],seed[1909],seed[3589],seed[3990],seed[2259],seed[552],seed[2137],seed[2417],seed[139],seed[1858],seed[30],seed[3379],seed[3909],seed[3353],seed[3661],seed[919],seed[314],seed[3255],seed[93],seed[94],seed[2263],seed[2439],seed[3225],seed[1363],seed[3783],seed[458],seed[2762],seed[1131],seed[1389],seed[2313],seed[310],seed[1851],seed[3637],seed[3126],seed[2628],seed[2155],seed[3808],seed[37],seed[3673],seed[3633],seed[3054],seed[2418],seed[841],seed[3668],seed[1355],seed[1515],seed[3039],seed[1714],seed[3960],seed[2593],seed[912],seed[1330],seed[3085],seed[1428],seed[409],seed[403],seed[915],seed[1267],seed[1904],seed[2824],seed[1050],seed[3655],seed[1784],seed[671],seed[2688],seed[3653],seed[3350],seed[3020],seed[2304],seed[844],seed[466],seed[3271],seed[206],seed[1846],seed[1077],seed[3935],seed[3779],seed[216],seed[40],seed[753],seed[622],seed[2190],seed[2332],seed[495],seed[1613],seed[735],seed[2208],seed[2774],seed[513],seed[1457],seed[3755],seed[977],seed[3123],seed[3538],seed[2614],seed[1900],seed[1703],seed[3967],seed[1451],seed[1265],seed[3798],seed[3660],seed[1029],seed[2710],seed[1149],seed[90],seed[2298],seed[3687],seed[3437],seed[2978],seed[2733],seed[1744],seed[3034],seed[280],seed[1864],seed[1512],seed[547],seed[3821],seed[99],seed[429],seed[2276],seed[1524],seed[1233],seed[1910],seed[3836],seed[3321],seed[1685],seed[1358],seed[3665],seed[1229],seed[3143],seed[2300],seed[3068],seed[1550],seed[1554],seed[2973],seed[3675],seed[2013],seed[1156],seed[2977],seed[2649],seed[1070],seed[3807],seed[2127],seed[284],seed[2475],seed[2696],seed[1508],seed[1469],seed[3438],seed[879],seed[2039],seed[366],seed[3723],seed[3997],seed[1540],seed[2136],seed[3406],seed[1388],seed[2491],seed[718],seed[3852],seed[1346],seed[3793],seed[831],seed[3331],seed[4002],seed[2838],seed[1083],seed[1939],seed[266],seed[3280],seed[106],seed[2312],seed[921],seed[2914],seed[956],seed[2296],seed[1255],seed[1867],seed[159],seed[937],seed[1545],seed[1810],seed[2187],seed[3448],seed[3885],seed[2207],seed[3879],seed[3847],seed[3943],seed[2324],seed[156],seed[1935],seed[2885],seed[3163],seed[2656],seed[2053],seed[2754],seed[854],seed[2396],seed[3443],seed[1391],seed[700],seed[3840],seed[1300],seed[853],seed[2171],seed[1422],seed[3611],seed[567],seed[2279],seed[1151],seed[1397],seed[3299],seed[2969],seed[1101],seed[907],seed[1369],seed[3302],seed[3801],seed[4080],seed[2815],seed[245],seed[1994],seed[2178],seed[2290],seed[3305],seed[1636],seed[1406],seed[2833],seed[2206],seed[1729],seed[4022],seed[2120],seed[3073],seed[2359],seed[866],seed[872],seed[2242],seed[684],seed[2745],seed[2703],seed[2956],seed[336],seed[1152],seed[3359],seed[2225],seed[2717],seed[766],seed[2452],seed[3995],seed[2151],seed[625],seed[3714],seed[1028],seed[3510],seed[278],seed[337],seed[3101],seed[4051],seed[1354],seed[2125],seed[431],seed[1412],seed[1787],seed[1199],seed[3874],seed[902],seed[2031],seed[2706],seed[1739],seed[2636],seed[2830],seed[2915],seed[3866],seed[2886],seed[721],seed[3659],seed[1294],seed[2468],seed[60],seed[1941],seed[235],seed[1244],seed[430],seed[2320],seed[2911],seed[319],seed[2965],seed[1332],seed[1668],seed[427],seed[1745],seed[2443],seed[604],seed[3129],seed[131],seed[2846],seed[2461],seed[1249],seed[2671],seed[1026],seed[258],seed[926],seed[1754],seed[3098],seed[1450],seed[50],seed[3449],seed[470],seed[1308],seed[2580],seed[1390],seed[170],seed[2597],seed[3692],seed[2801],seed[1727],seed[2613],seed[1023],seed[3062],seed[548],seed[2980],seed[351],seed[3566],seed[2212],seed[1110],seed[3090],seed[3501],seed[2749],seed[2447],seed[3499],seed[538],seed[2596],seed[2221],seed[808],seed[1608],seed[315],seed[3391],seed[3514],seed[2507],seed[2623],seed[3077],seed[3374],seed[1171],seed[1930],seed[4074],seed[1107],seed[2528],seed[3992],seed[3214],seed[393],seed[675],seed[3013],seed[594],seed[1018],seed[3833],seed[3677],seed[694],seed[1282],seed[1559],seed[2912],seed[3898],seed[4081],seed[2142],seed[2926],seed[693]}; 

//    end
    
    bsc bsc1(
        .clk(clk),
        .reset(reset),
        .seed({seed[1227],seed[2508],seed[1106],seed[543],seed[3292],seed[2432],seed[1097],seed[2437],seed[1154],seed[1644],seed[3327],seed[1620],seed[25],seed[1404],seed[2426],seed[1993],seed[463],seed[2638],seed[2804],seed[671],seed[927],seed[3516],seed[54],seed[7],seed[859],seed[648],seed[2616],seed[2593],seed[2880],seed[3772],seed[1755],seed[2394],seed[2021],seed[2525],seed[2233],seed[2965],seed[2323],seed[3719],seed[2167],seed[143],seed[1652],seed[990],seed[1495],seed[1220],seed[75],seed[2570],seed[202],seed[2014],seed[3864],seed[3013],seed[3214],seed[1998],seed[2296],seed[532],seed[523],seed[379],seed[3116],seed[1668],seed[1746],seed[695],seed[490],seed[3887],seed[3315],seed[2571],seed[3671],seed[3740],seed[2254],seed[1735],seed[1113],seed[2645],seed[1301],seed[23],seed[460],seed[253],seed[186],seed[3471],seed[3979],seed[893],seed[3350],seed[3570],seed[2642],seed[4056],seed[1233],seed[2791],seed[3421],seed[913],seed[2294],seed[158],seed[3794],seed[2895],seed[3591],seed[3764],seed[779],seed[1364],seed[4026],seed[3910],seed[3991],seed[218],seed[541],seed[1198],seed[3127],seed[1088],seed[670],seed[3707],seed[4086],seed[1875],seed[1325],seed[144],seed[2757],seed[113],seed[4054],seed[3607],seed[1509],seed[3282],seed[2382],seed[1419],seed[2983],seed[2482],seed[185],seed[1247],seed[2255],seed[1833],seed[1855],seed[615],seed[1557],seed[896],seed[3766],seed[1276],seed[2594],seed[562],seed[1929],seed[3807],seed[3852],seed[2524],seed[3552],seed[832],seed[3551],seed[2654],seed[940],seed[678],seed[2991],seed[276],seed[1067],seed[833],seed[1210],seed[3657],seed[888],seed[2945],seed[427],seed[3658],seed[3654],seed[3232],seed[898],seed[3435],seed[3888],seed[593],seed[518],seed[433],seed[3799],seed[660],seed[2690],seed[3099],seed[2583],seed[3792],seed[135],seed[169],seed[3999],seed[1902],seed[3021],seed[472],seed[1409],seed[3870],seed[1654],seed[3428],seed[181],seed[2313],seed[1188],seed[3086],seed[3128],seed[3094],seed[596],seed[232],seed[209],seed[3803],seed[3755],seed[2155],seed[3411],seed[2126],seed[1085],seed[2700],seed[2089],seed[2454],seed[340],seed[2213],seed[105],seed[3412],seed[2780],seed[96],seed[3083],seed[3381],seed[3631],seed[2451],seed[3301],seed[1141],seed[4042],seed[2103],seed[1104],seed[2678],seed[1546],seed[3082],seed[2116],seed[1624],seed[2694],seed[193],seed[2952],seed[3668],seed[2993],seed[2316],seed[3929],seed[2272],seed[821],seed[3268],seed[2201],seed[243],seed[1318],seed[1844],seed[617],seed[774],seed[819],seed[234],seed[2440],seed[439],seed[581],seed[527],seed[142],seed[1846],seed[2994],seed[1782],seed[134],seed[3366],seed[3946],seed[633],seed[2695],seed[1817],seed[569],seed[2207],seed[3394],seed[1921],seed[3944],seed[2276],seed[3811],seed[414],seed[509],seed[1870],seed[1759],seed[891],seed[422],seed[3859],seed[4],seed[466],seed[22],seed[822],seed[338],seed[3647],seed[3741],seed[2541],seed[2093],seed[1692],seed[2953],seed[3300],seed[2239],seed[1084],seed[1629],seed[2020],seed[1768],seed[2234],seed[3066],seed[2324],seed[281],seed[547],seed[634],seed[1825],seed[1293],seed[259],seed[520],seed[907],seed[1648],seed[97],seed[592],seed[2340],seed[1513],seed[174],seed[3734],seed[599],seed[2134],seed[2724],seed[1878],seed[2259],seed[3016],seed[3360],seed[1882],seed[291],seed[761],seed[428],seed[199],seed[628],seed[1715],seed[872],seed[1248],seed[2794],seed[407],seed[843],seed[2297],seed[3841],seed[3050],seed[279],seed[2310],seed[2264],seed[1723],seed[3184],seed[2876],seed[957],seed[3011],seed[842],seed[1436],seed[1559],seed[3438],seed[91],seed[2899],seed[2359],seed[180],seed[3558],seed[692],seed[258],seed[1476],seed[3917],seed[533],seed[2919],seed[3409],seed[1699],seed[1549],seed[1359],seed[1566],seed[2623],seed[3873],seed[3364],seed[2399],seed[1612],seed[3642],seed[3244],seed[392],seed[1901],seed[3967],seed[2818],seed[2946],seed[2352],seed[4091],seed[1679],seed[99],seed[1693],seed[1724],seed[2085],seed[1795],seed[398],seed[13],seed[231],seed[70],seed[3565],seed[1616],seed[2712],seed[487],seed[1398],seed[1353],seed[580],seed[4043],seed[1203],seed[489],seed[94],seed[840],seed[1176],seed[2607],seed[1029],seed[3156],seed[2873],seed[3203],seed[3983],seed[2446],seed[1414],seed[3957],seed[3447],seed[2867],seed[2223],seed[3492],seed[221],seed[1574],seed[2447],seed[3208],seed[3371],seed[29],seed[924],seed[3238],seed[133],seed[3161],seed[3387],seed[3950],seed[673],seed[1063],seed[3400],seed[2337],seed[3532],seed[697],seed[4068],seed[519],seed[1142],seed[1390],seed[1206],seed[1927],seed[3786],seed[4012],seed[557],seed[3334],seed[2245],seed[1886],seed[3056],seed[2069],seed[3134],seed[2145],seed[2746],seed[735],seed[2051],seed[2733],seed[81],seed[3789],seed[2332],seed[2626],seed[3470],seed[192],seed[227],seed[1773],seed[368],seed[1776],seed[1584],seed[920],seed[2606],seed[720],seed[3678],seed[1893],seed[3049],seed[1861],seed[1308],seed[2148],seed[828],seed[2967],seed[3320],seed[3069],seed[1483],seed[1672],seed[3927],seed[2424],seed[84],seed[3940],seed[3380],seed[1591],seed[2956],seed[892],seed[1857],seed[1610],seed[665],seed[1134],seed[986],seed[3439],seed[528],seed[1568],seed[2665],seed[3397],seed[900],seed[1479],seed[1722],seed[1767],seed[330],seed[1634],seed[1055],seed[3129],seed[3098],seed[1137],seed[1852],seed[1830],seed[2331],seed[3197],seed[3425],seed[2811],seed[3237],seed[3540],seed[383],seed[2191],seed[1018],seed[1793],seed[2681],seed[118],seed[3589],seed[3302],seed[1373],seed[2787],seed[2820],seed[4009],seed[2256],seed[352],seed[2403],seed[3923],seed[213],seed[559],seed[654],seed[1529],seed[3499],seed[4011],seed[1347],seed[4030],seed[3667],seed[2640],seed[984],seed[864],seed[579],seed[1717],seed[1528],seed[2909],seed[1785],seed[2949],seed[1482],seed[1384],seed[2793],seed[1408],seed[2664],seed[1897],seed[3026],seed[3939],seed[1499],seed[3139],seed[1473],seed[2462],seed[709],seed[1057],seed[611],seed[813],seed[1514],seed[3234],seed[3406],seed[2326],seed[1845],seed[1681],seed[2035],seed[2227],seed[3462],seed[384],seed[1890],seed[2445],seed[434],seed[3229],seed[2158],seed[825],seed[2796],seed[2822],seed[1311],seed[582],seed[1895],seed[1771],seed[3006],seed[2527],seed[139],seed[3575],seed[3079],seed[928],seed[2932],seed[851],seed[1952],seed[3716],seed[1205],seed[146],seed[385],seed[3791],seed[2143],seed[2305],seed[155],seed[469],seed[4064],seed[3919],seed[3801],seed[59],seed[788],seed[3963],seed[1928],seed[537],seed[3655],seed[542],seed[722],seed[3324],seed[2773],seed[2137],seed[3812],seed[223],seed[2784],seed[3624],seed[1996],seed[1385],seed[3926],seed[3760],seed[576],seed[1918],seed[2749],seed[393],seed[2769],seed[1268],seed[2772],seed[3019],seed[3553],seed[3456],seed[3988],seed[2529],seed[734],seed[2622],seed[1179],seed[3797],seed[2418],seed[175],seed[4093],seed[979],seed[1617],seed[1659],seed[1696],seed[3603],seed[1209],seed[3871],seed[1963],seed[2173],seed[2037],seed[1147],seed[2885],seed[103],seed[626],seed[3109],seed[3287],seed[2697],seed[2986],seed[3351],seed[1037],seed[2419],seed[436],seed[1231],seed[2829],seed[3155],seed[555],seed[3533],seed[2483],seed[1302],seed[3866],seed[1753],seed[1274],seed[1791],seed[621],seed[195],seed[587],seed[172],seed[3115],seed[1031],seed[3095],seed[3259],seed[170],seed[1720],seed[961],seed[1335],seed[1238],seed[1687],seed[1118],seed[3555],seed[3040],seed[2217],seed[3643],seed[4065],seed[3133],seed[1333],seed[3976],seed[1994],seed[306],seed[3293],seed[1326],seed[2547],seed[1619],seed[2591],seed[4057],seed[3121],seed[403],seed[3105],seed[3077],seed[72],seed[3557],seed[2628],seed[1809],seed[1168],seed[2834],seed[1937],seed[3452],seed[298],seed[2280],seed[2864],seed[3977],seed[3507],seed[2457],seed[1639],seed[246],seed[1818],seed[2602],seed[3503],seed[2067],seed[3743],seed[343],seed[1805],seed[2955],seed[2709],seed[753],seed[1425],seed[2146],seed[4017],seed[3189],seed[3487],seed[2325],seed[2110],seed[1540],seed[77],seed[3955],seed[1623],seed[3501],seed[3691],seed[2329],seed[3297],seed[3612],seed[2542],seed[4031],seed[1224],seed[3329],seed[3619],seed[566],seed[981],seed[1292],seed[121],seed[855],seed[2463],seed[4069],seed[3855],seed[2514],seed[2611],seed[3442],seed[723],seed[3798],seed[3395],seed[409],seed[1050],seed[2963],seed[1920],seed[2226],seed[3266],seed[1820],seed[2376],seed[3878],seed[1675],seed[1530],seed[2655],seed[442],seed[3032],seed[3247],seed[1502],seed[2502],seed[1150],seed[2300],seed[431],seed[3845],seed[3554],seed[1126],seed[3393],seed[1757],seed[2420],seed[2790],seed[1339],seed[3308],seed[705],seed[2806],seed[4052],seed[3168],seed[870],seed[3340],seed[1489],seed[1831],seed[4010],seed[3010],seed[3354],seed[2472],seed[1816],seed[3769],seed[2471],seed[1064],seed[110],seed[2357],seed[1909],seed[3055],seed[326],seed[3463],seed[295],seed[2507],seed[1307],seed[2936],seed[2042],seed[3973],seed[1058],seed[3166],seed[2598],seed[1714],seed[3593],seed[1321],seed[288],seed[2910],seed[539],seed[1520],seed[2208],seed[2004],seed[755],seed[1880],seed[680],seed[737],seed[3971],seed[3728],seed[2595],seed[2624],seed[2795],seed[3294],seed[3722],seed[1131],seed[553],seed[1285],seed[1907],seed[3724],seed[1941],seed[3897],seed[63],seed[3446],seed[701],seed[3997],seed[1556],seed[1636],seed[2985],seed[922],seed[650],seed[3260],seed[2676],seed[1152],seed[359],seed[2517],seed[1740],seed[353],seed[3020],seed[1627],seed[1704],seed[2520],seed[3907],seed[1649],seed[827],seed[1],seed[1609],seed[2609],seed[2816],seed[560],seed[3171],seed[2923],seed[1066],seed[1146],seed[911],seed[2815],seed[2738],seed[222],seed[1484],seed[1194],seed[3090],seed[2835],seed[2405],seed[1637],seed[770],seed[18],seed[1498],seed[1277],seed[767],seed[2311],seed[2767],seed[3683],seed[959],seed[205],seed[1362],seed[1047],seed[1828],seed[3521],seed[2629],seed[2212],seed[4040],seed[2088],seed[488],seed[885],seed[880],seed[980],seed[1580],seed[1647],seed[3935],seed[2590],seed[3508],seed[4087],seed[21],seed[3602],seed[196],seed[3932],seed[1433],seed[263],seed[563],seed[1177],seed[71],seed[3306],seed[1181],seed[3833],seed[3617],seed[2358],seed[1738],seed[3851],seed[292],seed[3921],seed[2289],seed[3249],seed[3213],seed[3087],seed[2801],seed[3182],seed[948],seed[405],seed[2027],seed[458],seed[1618],seed[1402],seed[4001],seed[610],seed[173],seed[1242],seed[1173],seed[3776],seed[1374],seed[2417],seed[1167],seed[3609],seed[3633],seed[3410],seed[974],seed[1917],seed[43],seed[2371],seed[1239],seed[2006],seed[3399],seed[2854],seed[3365],seed[3111],seed[2287],seed[381],seed[1216],seed[1544],seed[2355],seed[1581],seed[651],seed[3423],seed[416],seed[2937],seed[201],seed[93],seed[1615],seed[2969],seed[884],seed[3699],seed[1972],seed[2778],seed[2905],seed[3547],seed[2637],seed[2900],seed[2029],seed[3067],seed[3818],seed[3781],seed[2238],seed[3538],seed[661],seed[903],seed[3120],seed[797],seed[2510],seed[516],seed[3649],seed[360],seed[3909],seed[2001],seed[2277],seed[2040],seed[2762],seed[37],seed[3536],seed[1430],seed[3641],seed[1606],seed[1105],seed[2842],seed[1368],seed[4049],seed[2914],seed[1829],seed[423],seed[334],seed[117],seed[3383],seed[2858],seed[305],seed[4021],seed[3341],seed[3960],seed[841],seed[848],seed[3088],seed[1564],seed[679],seed[3338],seed[1860],seed[3986],seed[1748],seed[2187],seed[2667],seed[852],seed[3714],seed[507],seed[2597],seed[983],seed[3860],seed[3648],seed[130],seed[991],seed[2281],seed[1132],seed[2002],seed[255],seed[534],seed[20],seed[415],seed[3241],seed[1367],seed[1572],seed[718],seed[2828],seed[1447],seed[1360],seed[623],seed[3632],seed[3479],seed[787],seed[2916],seed[1645],seed[2630],seed[402],seed[2050],seed[1014],seed[785],seed[244],seed[2041],seed[2232],seed[2209],seed[491],seed[600],seed[782],seed[3936],seed[877],seed[760],seed[3461],seed[830],seed[3636],seed[1613],seed[1267],seed[1261],seed[2430],seed[696],seed[24],seed[260],seed[3690],seed[2499],seed[784],seed[2074],seed[741],seed[3024],seed[2468],seed[2601],seed[1330],seed[607],seed[3257],seed[3543],seed[283],seed[3753],seed[2887],seed[824],seed[1832],seed[2269],seed[2282],seed[2071],seed[3968],seed[742],seed[3071],seed[2157],seed[4006],seed[3969],seed[2713],seed[3408],seed[3686],seed[3842],seed[3065],seed[2328],seed[3829],seed[2200],seed[1211],seed[1357],seed[3018],seed[2861],seed[3003],seed[1734],seed[875],seed[3858],seed[1464],seed[1036],seed[1600],seed[2079],seed[40],seed[357],seed[3726],seed[4051],seed[3415],seed[1640],seed[3583],seed[4039],seed[1604],seed[814],seed[86],seed[3359],seed[854],seed[2843],seed[2911],seed[2260],seed[895],seed[2068],seed[1543],seed[2125],seed[2917],seed[2719],seed[646],seed[3270],seed[411],seed[1913],seed[938],seed[3494],seed[1579],seed[3809],seed[1096],seed[1287],seed[2752],seed[1388],seed[776],seed[1685],seed[3820],seed[1349],seed[1243],seed[2696],seed[2689],seed[1822],seed[2947],seed[3110],seed[881],seed[3418],seed[1214],seed[2186],seed[2774],seed[2679],seed[120],seed[2935],seed[3186],seed[2295],seed[1991],seed[3837],seed[2604],seed[1281],seed[2896],seed[1578],seed[733],seed[1790],seed[597],seed[3332],seed[1924],seed[1166],seed[4008],seed[3763],seed[1719],seed[1800],seed[2485],seed[2763],seed[2028],seed[1823],seed[479],seed[311],seed[603],seed[2240],seed[1508],seed[1827],seed[1742],seed[2782],seed[2384],seed[2727],seed[750],seed[3272],seed[1475],seed[3075],seed[1710],seed[3510],seed[441],seed[3876],seed[2686],seed[2308],seed[548],seed[1417],seed[2580],seed[769],seed[2532],seed[1535],seed[2109],seed[883],seed[3254],seed[1487],seed[2924],seed[128],seed[3243],seed[1560],seed[3444],seed[3250],seed[1836],seed[3277],seed[2195],seed[1080],seed[530],seed[1872],seed[3738],seed[627],seed[3634],seed[1076],seed[4025],seed[3422],seed[325],seed[1966],seed[3312],seed[1807],seed[2474],seed[1550],seed[3942],seed[1413],seed[2488],seed[745],seed[2996],seed[3046],seed[3718],seed[823],seed[585],seed[1752],seed[2734],seed[2184],seed[996],seed[1102],seed[4090],seed[2587],seed[3022],seed[3504],seed[2284],seed[2242],seed[1159],seed[3937],seed[987],seed[2862],seed[3733],seed[200],seed[3568],seed[1418],seed[3822],seed[1571],seed[1423],seed[3262],seed[480],seed[1949],seed[1303],seed[951],seed[282],seed[2064],seed[638],seed[2120],seed[2177],seed[4078],seed[1984],seed[316],seed[1358],seed[1389],seed[3037],seed[1381],seed[2721],seed[2731],seed[3154],seed[2224],seed[3588],seed[2891],seed[3629],seed[2452],seed[1300],seed[2768],seed[125],seed[64],seed[275],seed[3879],seed[3677],seed[3981],seed[3458],seed[3891],seed[1200],seed[2631],seed[3443],seed[52],seed[937],seed[304],seed[1053],seed[3496],seed[740],seed[2617],seed[2559],seed[80],seed[1938],seed[3062],seed[2270],seed[3373],seed[3747],seed[1153],seed[1183],seed[1437],seed[484],seed[588],seed[485],seed[4083],seed[2106],seed[2258],seed[2022],seed[1270],seed[656],seed[450],seed[1298],seed[529],seed[946],seed[167],seed[2391],seed[3271],seed[2298],seed[3356],seed[1077],seed[157],seed[2564],seed[2176],seed[3303],seed[2663],seed[1932],seed[3759],seed[3137],seed[0],seed[4070],seed[3],seed[449],seed[1427],seed[1667],seed[3468],seed[693],seed[2135],seed[2342],seed[207],seed[2413],seed[438],seed[1288],seed[3836],seed[2644],seed[1943],seed[3651],seed[2132],seed[1934],seed[2929],seed[274],seed[1232],seed[2379],seed[371],seed[1324],seed[1174],seed[2897],seed[1967],seed[2855],seed[1987],seed[3500],seed[3033],seed[1497],seed[3795],seed[2660],seed[1485],seed[2839],seed[2012],seed[3188],seed[3542],seed[2797],seed[2693],seed[3138],seed[3124],seed[2530],seed[2668],seed[1968],seed[1631],seed[932],seed[3093],seed[1969],seed[1350],seed[3278],seed[2998],seed[3349],seed[49],seed[214],seed[1850],seed[287],seed[1910],seed[3353],seed[1980],seed[2222],seed[2097],seed[210],seed[313],seed[2692],seed[224],seed[254],seed[3779],seed[1607],seed[3289],seed[3611],seed[3190],seed[2343],seed[3523],seed[690],seed[3970],seed[3497],seed[3073],seed[1130],seed[1702],seed[3592],seed[3493],seed[1611],seed[2557],seed[1678],seed[567],seed[2531],seed[2312],seed[290],seed[794],seed[982],seed[1810],seed[335],seed[1554],seed[2671],seed[796],seed[448],seed[1576],seed[2129],seed[3343],seed[2632],seed[2776],seed[577],seed[905],seed[3846],seed[4033],seed[2206],seed[3625],seed[3665],seed[150],seed[2330],seed[2438],seed[3585],seed[2095],seed[775],seed[3346],seed[3265],seed[406],seed[3347],seed[2718],seed[3159],seed[236],seed[916],seed[879],seed[3160],seed[1835],seed[1240],seed[1582],seed[1124],seed[3377],seed[2893],seed[2180],seed[219],seed[3001],seed[2183],seed[1575],seed[376],seed[2560],seed[1628],seed[3034],seed[1555],seed[2511],seed[1745],seed[1143],seed[3739],seed[417],seed[2056],seed[332],seed[3512],seed[554],seed[3045],seed[2883],seed[272],seed[2526],seed[4082],seed[358],seed[41],seed[3404],seed[2464],seed[2741],seed[4036],seed[2698],seed[453],seed[3749],seed[2049],seed[1761],seed[2759],seed[2901],seed[3267],seed[2725],seed[3630],seed[2387],seed[2026],seed[3194],seed[754],seed[2652],seed[2860],seed[3054],seed[1445],seed[3574],seed[3783],seed[1098],seed[267],seed[2516],seed[2119],seed[2484],seed[2107],seed[1521],seed[38],seed[866],seed[1492],seed[3269],seed[1320],seed[871],seed[389],seed[3273],seed[849],seed[2404],seed[2980],seed[296],seed[1565],seed[129],seed[2573],seed[16],seed[1283],seed[2635],seed[3118],seed[3616],seed[772],seed[2214],seed[853],seed[2024],seed[2651],seed[3736],seed[799],seed[3948],seed[2203],seed[2549],seed[319],seed[918],seed[252],seed[1586],seed[3370],seed[1252],seed[399],seed[437],seed[418],seed[1762],seed[2388],seed[771],seed[257],seed[2202],seed[3587],seed[1990],seed[1597],seed[2925],seed[1208],seed[3610],seed[3474],seed[1510],seed[3117],seed[978],seed[2467],seed[1642],seed[1093],seed[1501],seed[2052],seed[2448],seed[1455],seed[2096],seed[2370],seed[3869],seed[467],seed[3793],seed[3990],seed[2934],seed[1415],seed[2309],seed[3951],seed[3417],seed[3582],seed[882],seed[2592],seed[2179],seed[2962],seed[2237],seed[3815],seed[2892],seed[1522],seed[4095],seed[1770],seed[92],seed[1079],seed[455],seed[1854],seed[1100],seed[684],seed[2603],seed[1989],seed[2981],seed[2904],seed[2303],seed[934],seed[1392],seed[2301],seed[3255],seed[570],seed[1016],seed[1518],seed[1013],seed[1361],seed[2657],seed[3908],seed[1295],seed[2423],seed[2154],seed[1786],seed[1022],seed[2299],seed[668],seed[3701],seed[3856],seed[2216],seed[3051],seed[2168],seed[1342],seed[2252],seed[886],seed[3389],seed[1226],seed[1673],seed[3429],seed[909],seed[565],seed[2378],seed[944],seed[2572],seed[1467],seed[2821],seed[2008],seed[1784],seed[347],seed[369],seed[3502],seed[208],seed[3078],seed[1657],seed[1733],seed[2722],seed[61],seed[746],seed[2827],seed[1806],seed[837],seed[3113],seed[1906],seed[942],seed[874],seed[688],seed[2519],seed[1397],seed[1383],seed[3176],seed[3644],seed[3092],seed[3455],seed[2112],seed[2372],seed[1365],seed[2605],seed[3295],seed[2480],seed[3674],seed[1470],seed[2555],seed[85],seed[2044],seed[1936],seed[575],seed[3276],seed[459],seed[3027],seed[2427],seed[1382],seed[2845],seed[156],seed[598],seed[2927],seed[1466],seed[3253],seed[3645],seed[1780],seed[1663],seed[2215],seed[12],seed[618],seed[3918],seed[2118],seed[3322],seed[171],seed[1834],seed[3169],seed[56],seed[3445],seed[127],seed[3883],seed[2491],seed[2374],seed[1289],seed[2755],seed[8],seed[477],seed[413],seed[395],seed[624],seed[3985],seed[1265],seed[925],seed[154],seed[2055],seed[1869],seed[3828],seed[3331],seed[1935],seed[2979],seed[1481],seed[1655],seed[3806],seed[1751],seed[2381],seed[2278],seed[3219],seed[3752],seed[35],seed[3486],seed[613],seed[1337],seed[2128],seed[2354],seed[1109],seed[44],seed[1876],seed[998],seed[3344],seed[672],seed[4028],seed[2817],seed[2481],seed[1279],seed[1838],seed[27],seed[3785],seed[3835],seed[730],seed[1690],seed[309],seed[229],seed[2569],seed[2494],seed[1428],seed[3060],seed[3770],seed[230],seed[3639],seed[1898],seed[635],seed[114],seed[1212],seed[1336],seed[3978],seed[1983],seed[1169],seed[2477],seed[2150],seed[3672],seed[2080],seed[1553],seed[3717],seed[3142],seed[2961],seed[1879],seed[1658],seed[1865],seed[1905],seed[1450],seed[166],seed[2879],seed[710],seed[1567],seed[1583],seed[107],seed[1904],seed[1848],seed[2000],seed[2091],seed[3653],seed[2496],seed[2868],seed[2218],seed[2105],seed[1222],seed[1551],seed[2959],seed[3070],seed[969],seed[2551],seed[65],seed[3059],seed[106],seed[4059],seed[3945],seed[2992],seed[1074],seed[1766],seed[3413],seed[159],seed[2761],seed[1376],seed[2705],seed[3546],seed[2523],seed[1352],seed[2025],seed[1587],seed[4060],seed[57],seed[447],seed[34],seed[3029],seed[1725],seed[2383],seed[1033],seed[2841],seed[3482],seed[492],seed[3802],seed[2136],seed[3920],seed[3367],seed[2365],seed[3164],seed[3566],seed[3576],seed[2409],seed[2063],seed[1228],seed[2054],seed[67],seed[2625],seed[873],seed[3431],seed[2100],seed[3434],seed[3426],seed[3089],seed[867],seed[1071],seed[708],seed[985],seed[493],seed[2972],seed[504],seed[198],seed[1396],seed[3775],seed[2938],seed[1900],seed[1930],seed[2034],seed[3158],seed[3721],seed[876],seed[939],seed[564],seed[2647],seed[4007],seed[3746],seed[1032],seed[4089],seed[1442],seed[3601],seed[3025],seed[1314],seed[1923],seed[2402],seed[3572],seed[3831],seed[977],seed[3200],seed[2416],seed[1117],seed[1743],seed[2706],seed[540],seed[4050],seed[2369],seed[3378],seed[3626],seed[112],seed[1813],seed[1044],seed[248],seed[2567],seed[2509],seed[1674],seed[686],seed[691],seed[1970],seed[2292],seed[2009],seed[400],seed[496],seed[2826],seed[3005],seed[1925],seed[1887],seed[3898],seed[1729],seed[1812],seed[2246],seed[445],seed[2673],seed[2196],seed[1940],seed[950],seed[3074],seed[715],seed[4032],seed[2585],seed[1123],seed[3449],seed[2401],seed[2926],seed[857],seed[4023],seed[2730],seed[2831],seed[1056],seed[3141],seed[3012],seed[1371],seed[2521],seed[1908],seed[1682],seed[3192],seed[816],seed[3635],seed[2077],seed[2715],seed[926],seed[4081],seed[666],seed[2639],seed[2613],seed[3790],seed[3205],seed[747],seed[310],seed[1230],seed[4080],seed[3638],seed[2850],seed[674],seed[820],seed[1533],seed[1051],seed[3628],seed[4074],seed[1468],seed[153],seed[1421],seed[3526],seed[2265],seed[639],seed[3682],seed[1331],seed[1394],seed[1027],seed[2273],seed[2141],seed[62],seed[3152],seed[2373],seed[887],seed[2266],seed[869],seed[3949],seed[2497],seed[2030],seed[151],seed[2503],seed[2680],seed[126],seed[3467],seed[3044],seed[1236],seed[2500],seed[277],seed[131],seed[1244],seed[3476],seed[1792],seed[2353],seed[3505],seed[1922],seed[240],seed[1781],seed[2957],seed[268],seed[1511],seed[994],seed[2288],seed[2364],seed[3750],seed[2243],seed[2770],seed[2348],seed[2728],seed[804],seed[3123],seed[1278],seed[1662],seed[2389],seed[1945],seed[764],seed[3398],seed[3915],seed[3998],seed[815],seed[375],seed[3995],seed[1758],seed[3847],seed[3352],seed[1234],seed[3202],seed[464],seed[1112],seed[963],seed[2977],seed[1387],seed[3854],seed[3085],seed[1840],seed[3256],seed[3788],seed[2247],seed[2674],seed[2],seed[3311],seed[1976],seed[1665],seed[1814],seed[3709],seed[2575],seed[3135],seed[3737],seed[2964],seed[1115],seed[3615],seed[474],seed[2669],seed[2410],seed[3913],seed[675],seed[109],seed[1457],seed[526],seed[2837],seed[1175],seed[2533],seed[1089],seed[2720],seed[391],seed[3107],seed[1633],seed[2600],seed[846],seed[3531],seed[2553],seed[780],seed[2013],seed[3901],seed[3596],seed[2094],seed[1237],seed[2918],seed[2648],seed[3436],seed[3982],seed[2479],seed[719],seed[3966],seed[1120],seed[2807],seed[3843],seed[2138],seed[3172],seed[2833],seed[204],seed[2458],seed[1161],seed[410],seed[1561],seed[2274],seed[152],seed[2019],seed[1709],seed[3405],seed[3796],seed[3535],seed[707],seed[1266],seed[4075],seed[988],seed[1221],seed[1802],seed[1730],seed[972],seed[115],seed[1635],seed[2475],seed[2701],seed[2211],seed[1862],seed[1400],seed[3757],seed[952],seed[3206],seed[3685],seed[2059],seed[2115],seed[3207],seed[2775],seed[2251],seed[68],seed[2554],seed[3577],seed[315],seed[2812],seed[2033],seed[751],seed[1165],seed[3209],seed[2408],seed[706],seed[362],seed[2320],seed[233],seed[2263],seed[3545],seed[3830],seed[1946],seed[1107],seed[2318],seed[265],seed[2459],seed[2687],seed[3102],seed[3170],seed[2181],seed[2267],seed[2130],seed[1892],seed[2236],seed[714],seed[1703],seed[1839],seed[1046],seed[2546],seed[2261],seed[3893],seed[1092],seed[271],seed[968],seed[3882],seed[30],seed[187],seed[1191],seed[954],seed[1598],seed[1005],seed[1939],seed[1386],seed[2851],seed[1988],seed[3047],seed[4037],seed[3827],seed[264],seed[1125],seed[4055],seed[1081],seed[3149],seed[971],seed[235],seed[1821],seed[3711],seed[3742],seed[184],seed[1552],seed[1128],seed[3491],seed[1926],seed[478],seed[2073],seed[1114],seed[2166],seed[2087],seed[3038],seed[2920],seed[2053],seed[4016],seed[3961],seed[1355],seed[643],seed[2522],seed[162],seed[1344],seed[1465],seed[2174],seed[2058],seed[2810],seed[862],seed[1916],seed[73],seed[3787],seed[3941],seed[11],seed[3911],seed[2043],seed[1585],seed[2888],seed[1819],seed[1171],seed[2726],seed[2439],seed[1315],seed[3895],seed[732],seed[495],seed[1997],seed[468],seed[752],seed[2171],seed[1708],seed[834],seed[331],seed[1217],seed[1646],seed[237],seed[1894],seed[1195],seed[462],seed[440],seed[2205],seed[552],seed[676],seed[3586],seed[793],seed[404],seed[2066],seed[3178],seed[3224],seed[960],seed[1170],seed[486],seed[2487],seed[3824],seed[1779],seed[3490],seed[2661],seed[2133],seed[1193],seed[1023],seed[2544],seed[2341],seed[1182],seed[658],seed[1537],seed[2881],seed[501],seed[66],seed[2513],seed[572],seed[1853],seed[3825],seed[653],seed[344],seed[3333],seed[3361],seed[3745],seed[2460],seed[3126],seed[3725],seed[1269],seed[3488],seed[1688],seed[1446],seed[2743],seed[749],seed[931],seed[3153],seed[2380],seed[1933],seed[3305],seed[102],seed[1348],seed[2235],seed[3771],seed[3280],seed[685],seed[1004],seed[2345],seed[1877],seed[1593],seed[3345],seed[3286],seed[1866],seed[1769],seed[1680],seed[763],seed[583],seed[3618],seed[420],seed[2366],seed[2204],seed[1523],seed[1881],seed[818],seed[3661],seed[3225],seed[2377],seed[2562],seed[289],seed[901],seed[2436],seed[3459],seed[3692],seed[3336],seed[1496],seed[1975],seed[179],seed[3712],seed[1366],seed[1911],seed[3518],seed[910],seed[3903],seed[2675],seed[1178],seed[3506],seed[1884],seed[682],seed[861],seed[3804],seed[3106],seed[1042],seed[728],seed[3465],seed[1562],seed[783],seed[2906],seed[1889],seed[836],seed[1686],seed[1858],seed[2540],seed[2392],seed[168],seed[293],seed[3819],seed[124],seed[3198],seed[1622],seed[844],seed[2007],seed[574],seed[620],seed[312],seed[2866],seed[3868],seed[811],seed[285],seed[372],seed[2225],seed[2882],seed[2819],seed[206],seed[1160],seed[2321],seed[3328],seed[1189],seed[2688],seed[2160],seed[941],seed[1985],seed[713],seed[1316],seed[3778],seed[808],seed[947],seed[3663],seed[147],seed[299],seed[2646],seed[1641],seed[294],seed[3478],seed[1590],seed[3342],seed[3623],seed[2621],seed[203],seed[3177],seed[88],seed[3689],seed[1973],seed[2199],seed[83],seed[4048],seed[3666],seed[3974],seed[3758],seed[2147],seed[777],seed[2090],seed[87],seed[1999],seed[663],seed[1246],seed[3727],seed[1062],seed[3520],seed[1713],seed[546],seed[374],seed[2633],seed[95],seed[1258],seed[894],seed[531],seed[3240],seed[2933],seed[1558],seed[100],seed[738],seed[3890],seed[602],seed[1180],seed[863],seed[970],seed[995],seed[1328],seed[2849],seed[2518],seed[1532],seed[3777],seed[1393],seed[2886],seed[2931],seed[2528],seed[3605],seed[3464],seed[3368],seed[3865],seed[538],seed[2512],seed[242],seed[3627],seed[1977],seed[3599],seed[2968],seed[161],seed[2290],seed[3580],seed[3216],seed[2971],seed[3402],seed[2162],seed[339],seed[1327],seed[3009],seed[1006],seed[3433],seed[3480],seed[1515],seed[4035],seed[2250],seed[3119],seed[2036],seed[1135],seed[2262],seed[2997],seed[2871],seed[1506],seed[3684],seed[182],seed[1061],seed[1797],seed[1486],seed[1136],seed[1015],seed[3659],seed[1341],seed[2574],seed[917],seed[2017],seed[9],seed[3251],seed[2170],seed[2057],seed[2443],seed[976],seed[2065],seed[1354],seed[1488],seed[3881],seed[845],seed[2039],seed[4015],seed[1859],seed[3773],seed[2102],seed[790],seed[524],seed[1025],seed[3076],seed[657],seed[3573],seed[997],seed[662],seed[1249],seed[3372],seed[435],seed[3097],seed[4047],seed[3556],seed[3309],seed[3813],seed[3694],seed[498],seed[3475],seed[3703],seed[1070],seed[1461],seed[1313],seed[1747],seed[1363],seed[3756],seed[386],seed[1961],seed[2407],seed[55],seed[2543],seed[739],seed[2393],seed[3840],seed[3637],seed[3564],seed[3730],seed[3140],seed[457],seed[256],seed[878],seed[625],seed[1028],seed[426],seed[2390],seed[999],seed[1286],seed[4071],seed[266],seed[3762],seed[3386],seed[380],seed[2535],seed[4077],seed[2178],seed[1040],seed[1202],seed[2588],seed[3191],seed[3581],seed[432],seed[545],seed[3318],seed[1503],seed[42],seed[1538],seed[2942],seed[1111],seed[2275],seed[1841],seed[2536],seed[3039],seed[2349],seed[101],seed[1103],seed[2940],seed[1660],seed[1312],seed[3004],seed[1605],seed[1694],seed[2060],seed[1959],seed[3290],seed[3590],seed[4002],seed[378],seed[317],seed[1643],seed[1405],seed[3880],seed[1356],seed[2156],seed[792],seed[3385],seed[2414],seed[1737],seed[3875],seed[3245],seed[3002],seed[614],seed[1669],seed[2185],seed[664],seed[558],seed[2677],seed[2431],seed[2608],seed[3849],seed[388],seed[1219],seed[2197],seed[3906],seed[3650],seed[2771],seed[2872],seed[3008],seed[3220],seed[762],seed[2825],seed[2003],seed[1676],seed[966],seed[2283],seed[1653],seed[3992],seed[341],seed[1625],seed[3481],seed[3183],seed[1749],seed[1218],seed[2104],seed[2747],seed[226],seed[4022],seed[1151],seed[1420],seed[2515],seed[3548],seed[3130],seed[3472],seed[4067],seed[3028],seed[3157],seed[2465],seed[51],seed[2078],seed[3620],seed[1310],seed[262],seed[1213],seed[2489],seed[2221],seed[2534],seed[3239],seed[3041],seed[3702],seed[1948],seed[342],seed[3061],seed[3030],seed[2010],seed[2788],seed[3321],seed[1411],seed[2350],seed[3103],seed[2783],seed[1078],seed[3457],seed[145],seed[3621],seed[616],seed[3180],seed[801],seed[2941],seed[1500],seed[3867],seed[3357],seed[3930],seed[1888],seed[322],seed[3477],seed[1319],seed[3195],seed[3081],seed[1626],seed[2113],seed[1808],seed[3780],seed[515],seed[3989],seed[647],seed[2466],seed[1458],seed[681],seed[3544],seed[550],seed[1577],seed[1589],seed[3165],seed[640],seed[2492],seed[2307],seed[4094],seed[953],seed[2684],seed[3122],seed[2636],seed[2153],seed[1187],seed[301],seed[1144],seed[2982],seed[1451],seed[3765],seed[2578],seed[1986],seed[2375],seed[280],seed[1121],seed[3975],seed[1273],seed[3104],seed[3928],seed[1684],seed[1380],seed[1811],seed[3705],seed[3330],seed[2428],seed[2581],seed[286],seed[1329],seed[2476],seed[3136],seed[2903],seed[3511],seed[3227],seed[703],seed[506],seed[1020],seed[2970],seed[250],seed[3774],seed[2351],seed[4005],seed[3108],seed[3660],seed[1095],seed[3844],seed[908],seed[2915],seed[2188],seed[2398],seed[2599],seed[1596],seed[328],seed[2169],seed[183],seed[3515],seed[3838],seed[1525],seed[2803],seed[2857],seed[4024],seed[3187],seed[3035],seed[1343],seed[4034],seed[212],seed[1410],seed[1296],seed[3112],seed[2335],seed[1192],seed[3369],seed[3744],seed[2415],seed[1241],seed[2228],seed[3222],seed[3114],seed[689],seed[3933],seed[470],seed[1148],seed[511],seed[586],seed[46],seed[1001],seed[631],seed[3162],seed[669],seed[1003],seed[2442],seed[2190],seed[3023],seed[3231],seed[261],seed[2083],seed[17],seed[3048],seed[812],seed[136],seed[3708],seed[1406],seed[390],seed[3877],seed[3823],seed[2653],seed[270],seed[958],seed[936],seed[1116],seed[2789],seed[2754],seed[1372],seed[164],seed[1264],seed[2385],seed[3952],seed[1731],seed[1978],seed[636],seed[397],seed[3640],seed[2944],seed[3199],seed[956],seed[1545],seed[1815],seed[1601],seed[3221],seed[2456],seed[1172],seed[1958],seed[3317],seed[2045],seed[1891],seed[2750],seed[3235],seed[3956],seed[39],seed[765],seed[2662],seed[2123],seed[1334],seed[45],seed[3695],seed[2271],seed[889],seed[3242],seed[2194],seed[3167],seed[1531],seed[2046],seed[1536],seed[3698],seed[2302],seed[3466],seed[3550],seed[2362],seed[2220],seed[1783],seed[249],seed[1962],seed[278],seed[930],seed[1035],seed[791],seed[929],seed[1796],seed[3248],seed[2966],seed[2634],seed[2455],seed[795],seed[2785],seed[3934],seed[1290],seed[1011],seed[1491],seed[3598],seed[2411],seed[425],seed[1275],seed[1008],seed[1801],seed[228],seed[284],seed[1774],seed[1251],seed[1305],seed[655],seed[1956],seed[2098],seed[1856],seed[2360],seed[4092],seed[3424],seed[2805],seed[1914],seed[3326],seed[2659],seed[4062],seed[1689],seed[1434],seed[412],seed[2576],seed[2586],seed[1664],seed[1030],seed[1982],seed[3145],seed[3100],seed[935],seed[622],seed[2751],seed[3440],seed[2877],seed[517],seed[419],seed[1896],seed[2610],seed[1379],seed[1260],seed[3484],seed[3007],seed[3959],seed[333],seed[2975],seed[3258],seed[1992],seed[1651],seed[1505],seed[497],seed[2612],seed[3862],seed[430],seed[2347],seed[1204],seed[3291],seed[3816],seed[1493],seed[141],seed[3212],seed[2429],seed[1947],seed[2682],seed[3376],seed[3509],seed[2386],seed[989],seed[321],seed[3965],seed[2809],seed[1794],seed[1199],seed[2737],seed[2939],seed[3335],seed[858],seed[1683],seed[778],seed[3252],seed[429],seed[1775],seed[768],seed[499],seed[3850],seed[3469],seed[2368],seed[632],seed[2249],seed[3652],seed[3519],seed[2334],seed[3285],seed[3473],seed[1534],seed[3375],seed[727],seed[1422],seed[111],seed[1843],seed[1122],seed[1424],seed[3264],seed[1750],seed[1441],seed[3441],seed[211],seed[2708],seed[3432],seed[2493],seed[3163],seed[1431],seed[1304],seed[1599],seed[759],seed[1705],seed[3430],seed[2930],seed[2649],seed[336],seed[2253],seed[590],seed[1739],seed[1259],seed[2824],seed[2047],seed[2650],seed[3800],seed[1282],seed[595],seed[2229],seed[810],seed[2890],seed[2434],seed[216],seed[1547],seed[2241],seed[475],seed[2257],seed[3233],seed[856],seed[2765],seed[494],seed[1912],seed[217],seed[1082],seed[2707],seed[1885],seed[1592],seed[2490],seed[1412],seed[2139],seed[965],seed[630],seed[3358],seed[1054],seed[245],seed[955],seed[451],seed[2954],seed[933],seed[4004],seed[2075],seed[4045],seed[149],seed[2683],seed[4053],seed[138],seed[2732],seed[2753],seed[1019],seed[4066],seed[644],seed[2248],seed[3052],seed[3896],seed[3147],seed[1697],seed[850],seed[297],seed[505],seed[60],seed[1127],seed[3569],seed[2672],seed[123],seed[1873],seed[2563],seed[2846],seed[4019],seed[839],seed[2461],seed[1691],seed[2444],seed[1711],seed[364],seed[373],seed[2950],seed[805],seed[3522],seed[2566],seed[1073],seed[1463],seed[1229],seed[1297],seed[2161],seed[1798],seed[4029],seed[3885],seed[1516],seed[1548],seed[3263],seed[606],seed[716],seed[3323],seed[3597],seed[3304],seed[251],seed[1614],seed[510],seed[2396],seed[3784],seed[1045],seed[1744],seed[3578],seed[1700],seed[2018],seed[3513],seed[4085],seed[90],seed[215],seed[365],seed[1039],seed[2121],seed[3299],seed[694],seed[2814],seed[2922],seed[1569],seed[1157],seed[1375],seed[773],seed[302],seed[2076],seed[1416],seed[2306],seed[3720],seed[1453],seed[2756],seed[1284],seed[1101],seed[3015],seed[140],seed[1849],seed[1460],seed[2114],seed[354],seed[1804],seed[377],seed[1155],seed[1507],seed[2230],seed[2397],seed[744],seed[3972],seed[2545],seed[1017],seed[1322],seed[3916],seed[659],seed[351],seed[104],seed[923],seed[3296],seed[4061],seed[2548],seed[2449],seed[137],seed[79],seed[1477],seed[798],seed[1524],seed[2092],seed[1608],seed[1378],seed[1443],seed[1826],seed[806],seed[1474],seed[2840],seed[3872],seed[452],seed[3731],seed[1254],seed[3680],seed[1778],seed[2422],seed[178],seed[641],seed[3058],seed[1440],seed[2870],seed[2131],seed[3420],seed[2579],seed[1139],seed[160],seed[1235],seed[3863],seed[2987],seed[712],seed[1883],seed[1456],seed[3261],seed[1971],seed[503],seed[4018],seed[3924],seed[3283],seed[561],seed[700],seed[3528],seed[2061],seed[1438],seed[2501],seed[241],seed[163],seed[1021],seed[3042],seed[1957],seed[2011],seed[3889],seed[2802],seed[1129],seed[2865],seed[2005],seed[1432],seed[3173],seed[2584],seed[3448],seed[2400],seed[789],seed[2670],seed[1317],seed[2568],seed[1162],seed[2286],seed[1294],seed[3943],seed[2729],seed[1863],seed[318],seed[2777],seed[1995],seed[2140],seed[1000],seed[2099],seed[1494],seed[2117],seed[2656],seed[786],seed[3101],seed[58],seed[2643],seed[2304],seed[3451],seed[36],seed[573],seed[3853],seed[1186],seed[3848],seed[3808],seed[1698],seed[3319],seed[2702],seed[3414],seed[3595],seed[1760],seed[2908],seed[4038],seed[3150],seed[2101],seed[2976],seed[3902],seed[2620],seed[3839],seed[1526],seed[2874],seed[2565],seed[3091],seed[482],seed[1185],seed[1837],seed[758],seed[2210],seed[1009],seed[1256],seed[781],seed[1280],seed[3325],seed[483],seed[1306],seed[4063],seed[3193],seed[1728],seed[3210],seed[571],seed[2658],seed[108],seed[2023],seed[3175],seed[645],seed[2948],seed[1184],seed[2974],seed[1944],seed[1435],seed[1931],seed[3401],seed[3754],seed[3805],seed[3761],seed[1541],seed[500],seed[1542],seed[2989],seed[591],seed[717],seed[2425],seed[4088],seed[3211],seed[1024],seed[421],seed[1661],seed[2710],seed[348],seed[3392],seed[612],seed[1951],seed[2627],seed[15],seed[1701],seed[3904],seed[2760],seed[2863],seed[1403],seed[1954],seed[704],seed[3579],seed[2291],seed[3673],seed[2015],seed[3886],seed[1156],seed[3382],seed[2641],seed[2764],seed[803],seed[3017],seed[1038],seed[3922],seed[3810],seed[461],seed[3179],seed[629],seed[589],seed[1223],seed[2149],seed[2781],seed[2152],seed[3832],seed[2082],seed[1452],seed[2907],seed[1656],seed[943],seed[3964],seed[1650],seed[446],seed[1824],seed[1588],seed[197],seed[1158],seed[3549],seed[2958],seed[512],seed[3228],seed[3236],seed[1960],seed[4020],seed[350],seed[2084],seed[1094],seed[1842],seed[829],seed[1964],seed[189],seed[3316],seed[1049],seed[3348],seed[1573],seed[619],seed[3606],seed[2293],seed[188],seed[1718],seed[2704],seed[3246],seed[3767],seed[3185],seed[382],seed[1765],seed[1271],seed[3201],seed[1108],seed[3064],seed[2193],seed[2798],seed[346],seed[1149],seed[973],seed[3676],seed[2314],seed[2470],seed[1272],seed[2716],seed[2847],seed[2577],seed[122],seed[33],seed[992],seed[3925],seed[1263],seed[1764],seed[525],seed[2744],seed[3388],seed[3374],seed[2219],seed[2124],seed[807],seed[247],seed[1763],seed[1091],seed[1519],seed[471],seed[702],seed[3892],seed[3947],seed[4046],seed[3537],seed[2538],seed[2766],seed[116],seed[1490],seed[3693],seed[1346],seed[78],seed[2995],seed[3530],seed[2031],seed[2736],seed[2127],seed[2315],seed[239],seed[3284],seed[502],seed[82],seed[3529],seed[176],seed[3748],seed[1083],seed[1439],seed[2182],seed[677],seed[838],seed[2159],seed[320],seed[3732],seed[1979],seed[1351],seed[3391],seed[3226],seed[551],seed[1340],seed[1632],seed[2361],seed[4044],seed[3313],seed[2421],seed[2504],seed[2327],seed[4079],seed[2441],seed[667],seed[3407],seed[3223],seed[2469],seed[363],seed[225],seed[3144],seed[835],seed[1090],seed[3700],seed[897],seed[3485],seed[1732],seed[2478],seed[3931],seed[1338],seed[2875],seed[3681],seed[1754],seed[2558],seed[1867],seed[1868],seed[3217],seed[3527],seed[2192],seed[324],seed[1727],seed[2723],seed[2832],seed[1196],seed[2990],seed[14],seed[1471],seed[2363],seed[3604],seed[2943],seed[2884],seed[3218],seed[860],seed[1060],seed[890],seed[2198],seed[26],seed[3600],seed[1010],seed[642],seed[1245],seed[1512],seed[2748],seed[4041],seed[4000],seed[1448],seed[1864],seed[3704],seed[6],seed[736],seed[3768],seed[711],seed[2108],seed[3396],seed[2921],seed[2506],seed[3403],seed[2086],seed[2336],seed[1190],seed[1981],seed[2435],seed[3125],seed[1119],seed[2703],seed[1472],seed[3814],seed[2163],seed[1459],seed[3987],seed[3524],seed[1429],seed[513],seed[2984],seed[1915],seed[47],seed[1603],seed[1594],seed[1145],seed[3498],seed[1087],seed[238],seed[3307],seed[424],seed[1670],seed[3894],seed[3416],seed[3584],seed[2164],seed[2836],seed[1695],seed[687],seed[3697],seed[2231],seed[2319],seed[2735],seed[3562],seed[465],seed[721],seed[69],seed[4072],seed[1323],seed[1630],seed[3900],seed[349],seed[3080],seed[2848],seed[847],seed[2172],seed[3131],seed[76],seed[3274],seed[3914],seed[98],seed[1257],seed[1426],seed[3817],seed[307],seed[766],seed[2618],seed[556],seed[3298],seed[1068],seed[19],seed[699],seed[2473],seed[2691],seed[2539],seed[1974],seed[148],seed[2016],seed[2338],seed[481],seed[3337],seed[1164],seed[1207],seed[3450],seed[303],seed[2556],seed[2537],seed[3072],seed[132],seed[865],seed[366],seed[902],seed[1369],seed[3594],seed[726],seed[3646],seed[2268],seed[1262],seed[2285],seed[269],seed[1851],seed[1138],seed[1401],seed[2142],seed[396],seed[1741],seed[3560],seed[1539],seed[367],seed[1299],seed[308],seed[817],seed[594],seed[1919],seed[1803],seed[3096],seed[1075],seed[2070],seed[3857],seed[2685],seed[3279],seed[2356],seed[3670],seed[2999],seed[1012],seed[2878],seed[3561],seed[975],seed[605],seed[1602],seed[3419],seed[3196],seed[89],seed[3899],seed[300],seed[3437],seed[1517],seed[3390],seed[1621],seed[355],seed[3706],seed[637],seed[1570],seed[2792],seed[3355],seed[2779],seed[370],seed[454],seed[53],seed[3363],seed[3204],seed[3427],seed[725],seed[3483],seed[1777],seed[2550],seed[2714],seed[2902],seed[2889],seed[1048],seed[2322],seed[1871],seed[1955],seed[2869],seed[2853],seed[2740],seed[3362],seed[3514],seed[2800],seed[1953],seed[1950],seed[1215],seed[906],seed[609],seed[3559],seed[456],seed[3614],seed[3068],seed[2898],seed[649],seed[3132],seed[964],seed[3053],seed[1899],seed[220],seed[2582],seed[508],seed[1309],seed[2838],seed[535],seed[2615],seed[329],seed[177],seed[1395],seed[2739],seed[3057],seed[119],seed[1007],seed[522],seed[3912],seed[2038],seed[1716],seed[3735],seed[3310],seed[2823],seed[756],seed[4027],seed[2367],seed[4084],seed[1026],seed[473],seed[809],seed[3000],seed[2333],seed[1462],seed[1399],seed[1480],seed[1903],seed[1407],seed[993],seed[337],seed[962],seed[2081],seed[3148],seed[1069],seed[802],seed[2619],seed[2589],seed[2856],seed[2433],seed[2928],seed[2813],seed[2175],seed[1706],seed[1391],seed[743],seed[327],seed[1345],seed[1677],seed[2032],seed[394],seed[3994],seed[3861],seed[4014],seed[1197],seed[899],seed[3453],seed[1332],seed[1787],seed[2758],seed[3275],seed[3723],seed[3143],seed[1250],seed[194],seed[4058],seed[3884],seed[28],seed[1527],seed[1253],seed[3339],seed[904],seed[2978],seed[3288],seed[1707],seed[2852],seed[1736],seed[2317],seed[3151],seed[3874],seed[514],seed[3954],seed[1726],seed[1942],seed[3826],seed[361],seed[2165],seed[1377],seed[345],seed[2894],seed[1454],seed[3181],seed[1002],seed[831],seed[3710],seed[1444],seed[1788],seed[3454],seed[2244],seed[826],seed[3517],seed[1201],seed[757],seed[3938],seed[1059],seed[3962],seed[2111],seed[50],seed[1086],seed[3669],seed[2912],seed[3541],seed[2859],seed[568],seed[2450],seed[2453],seed[915],seed[731],seed[1140],seed[2951],seed[444],seed[921],seed[945],seed[1469],seed[2913],seed[10],seed[2122],seed[2699],seed[1789],seed[3953],seed[578],seed[1041],seed[356],seed[967],seed[3993],seed[2614],seed[2666],seed[800],seed[2072],seed[2062],seed[1504],seed[1034],seed[2344],seed[2742],seed[165],seed[2745],seed[3539],seed[1595],seed[3613],seed[608],seed[1133],seed[1638],seed[1072],seed[2498],seed[32],seed[1666],seed[521],seed[1478],seed[1110],seed[2988],seed[3782],seed[3687],seed[2412],seed[604],seed[1052],seed[1756],seed[3146],seed[314],seed[3063],seed[2048],seed[3043],seed[3821],seed[2596],seed[4073],seed[912],seed[443],seed[536],seed[3905],seed[3215],seed[191],seed[2561],seed[2189],seed[190],seed[3656],seed[2406],seed[2346],seed[3563],seed[3834],seed[3230],seed[2717],seed[2973],seed[4013],seed[2339],seed[1370],seed[3958],seed[2144],seed[868],seed[1291],seed[3489],seed[74],seed[1772],seed[2279],seed[5],seed[4076],seed[584],seed[2552],seed[3664],seed[2395],seed[2505],seed[1563],seed[31],seed[3379],seed[3036],seed[2960],seed[914],seed[1099],seed[3014],seed[1965],seed[3713],seed[729],seed[3622],seed[3314],seed[748],seed[1449],seed[3384],seed[2151],seed[3495],seed[2486],seed[2830],seed[1721],seed[3996],seed[3675],seed[3696],seed[3031],seed[1043],seed[3567],seed[3980],seed[1225],seed[1712],seed[4003],seed[1255],seed[3984],seed[3608],seed[1065],seed[724],seed[1799],seed[1874],seed[3084],seed[1847],seed[2786],seed[2844],seed[683],seed[3534],seed[949],seed[3688],seed[698],seed[2495],seed[3525],seed[3571],seed[3281],seed[476],seed[3715],seed[601],seed[919],seed[387],seed[2808],seed[2711],seed[323],seed[48],seed[549],seed[1163],seed[544],seed[3460],seed[1671],seed[3751],seed[273],seed[3174],seed[401],seed[3662],seed[408],seed[3679],seed[2799],seed[3729],seed[652]}),
        .cross_prob(cross_prob),
        .codeword(codeword1),
        .received(received1)
        );
    
    bsc bsc2(
        .clk(clk),
        .reset(reset),
        .seed({seed[3755],seed[988],seed[3960],seed[2859],seed[2044],seed[1829],seed[2116],seed[1015],seed[1573],seed[1704],seed[2775],seed[3485],seed[652],seed[3089],seed[3870],seed[2905],seed[697],seed[1077],seed[1635],seed[2457],seed[1786],seed[337],seed[2174],seed[101],seed[2450],seed[3605],seed[2850],seed[2035],seed[2159],seed[3982],seed[1114],seed[3291],seed[3289],seed[3535],seed[1626],seed[1554],seed[853],seed[748],seed[1319],seed[1394],seed[3878],seed[2749],seed[689],seed[129],seed[1527],seed[3544],seed[590],seed[1489],seed[3025],seed[3055],seed[187],seed[3351],seed[744],seed[814],seed[507],seed[1270],seed[2474],seed[2639],seed[2600],seed[1353],seed[2841],seed[598],seed[3751],seed[1558],seed[3747],seed[1323],seed[746],seed[1875],seed[2814],seed[800],seed[4054],seed[1390],seed[180],seed[3702],seed[1134],seed[1138],seed[761],seed[874],seed[3410],seed[3995],seed[3958],seed[416],seed[4061],seed[3700],seed[585],seed[1706],seed[2538],seed[733],seed[2874],seed[1736],seed[449],seed[985],seed[2307],seed[54],seed[1898],seed[712],seed[3431],seed[856],seed[150],seed[727],seed[1537],seed[774],seed[1305],seed[2867],seed[2722],seed[721],seed[2616],seed[1284],seed[2017],seed[1456],seed[68],seed[2106],seed[4089],seed[3593],seed[1686],seed[364],seed[208],seed[2570],seed[919],seed[1940],seed[3326],seed[1079],seed[880],seed[3484],seed[961],seed[3411],seed[2279],seed[495],seed[888],seed[1807],seed[3013],seed[2382],seed[1619],seed[2120],seed[1004],seed[1980],seed[2950],seed[1605],seed[297],seed[2322],seed[3518],seed[1989],seed[1910],seed[1580],seed[2014],seed[1225],seed[1974],seed[506],seed[1876],seed[3557],seed[3369],seed[3546],seed[1363],seed[3770],seed[4035],seed[2624],seed[2271],seed[3576],seed[3930],seed[665],seed[1239],seed[3395],seed[3111],seed[3365],seed[3635],seed[2986],seed[3421],seed[3831],seed[2376],seed[312],seed[1998],seed[1287],seed[3683],seed[1852],seed[1480],seed[661],seed[1691],seed[3618],seed[1006],seed[3667],seed[2261],seed[4030],seed[1497],seed[244],seed[340],seed[3904],seed[3820],seed[2419],seed[1911],seed[1777],seed[3743],seed[1314],seed[3956],seed[3312],seed[1016],seed[350],seed[1375],seed[1117],seed[3246],seed[3631],seed[2893],seed[1423],seed[3415],seed[2422],seed[39],seed[3465],seed[3414],seed[1279],seed[2223],seed[2292],seed[2621],seed[3451],seed[3556],seed[3693],seed[1013],seed[1962],seed[3745],seed[715],seed[618],seed[3496],seed[3974],seed[2987],seed[3838],seed[2999],seed[3200],seed[3052],seed[140],seed[1514],seed[1630],seed[2104],seed[351],seed[4057],seed[4060],seed[2585],seed[1106],seed[3458],seed[1121],seed[957],seed[3595],seed[3638],seed[2448],seed[964],seed[656],seed[1377],seed[1078],seed[863],seed[1740],seed[2804],seed[1281],seed[2820],seed[2612],seed[807],seed[1617],seed[3011],seed[1871],seed[1930],seed[1470],seed[2752],seed[3066],seed[3021],seed[1963],seed[3905],seed[3777],seed[2015],seed[605],seed[1830],seed[2598],seed[2653],seed[1792],seed[135],seed[2484],seed[829],seed[2695],seed[1419],seed[2383],seed[2206],seed[3876],seed[430],seed[182],seed[3252],seed[1739],seed[3007],seed[1929],seed[250],seed[1559],seed[1782],seed[367],seed[594],seed[2565],seed[1757],seed[629],seed[1781],seed[824],seed[3785],seed[3815],seed[3215],seed[846],seed[3714],seed[927],seed[305],seed[3146],seed[2561],seed[3071],seed[3599],seed[4049],seed[3880],seed[3294],seed[3726],seed[1943],seed[3076],seed[553],seed[3059],seed[1009],seed[2700],seed[510],seed[2034],seed[2471],seed[59],seed[3773],seed[2916],seed[959],seed[2493],seed[749],seed[3727],seed[418],seed[282],seed[546],seed[262],seed[3340],seed[96],seed[3711],seed[338],seed[2674],seed[2951],seed[539],seed[3148],seed[3017],seed[693],seed[3607],seed[429],seed[2808],seed[2053],seed[840],seed[3302],seed[1436],seed[1841],seed[1324],seed[986],seed[1112],seed[319],seed[138],seed[3429],seed[3695],seed[516],seed[3149],seed[3166],seed[2851],seed[706],seed[1195],seed[2529],seed[4083],seed[2932],seed[1049],seed[222],seed[384],seed[163],seed[2890],seed[2815],seed[969],seed[1799],seed[291],seed[3975],seed[2954],seed[1442],seed[2944],seed[34],seed[467],seed[3152],seed[3416],seed[3924],seed[531],seed[3268],seed[2679],seed[4062],seed[1250],seed[595],seed[675],seed[153],seed[1310],seed[2738],seed[3664],seed[2568],seed[315],seed[2154],seed[2233],seed[2756],seed[3676],seed[1627],seed[3879],seed[520],seed[3996],seed[3644],seed[236],seed[2992],seed[1027],seed[2998],seed[1298],seed[2548],seed[827],seed[1268],seed[1304],seed[1983],seed[869],seed[3571],seed[2761],seed[809],seed[2193],seed[69],seed[3792],seed[3186],seed[698],seed[3629],seed[2681],seed[162],seed[3944],seed[1482],seed[3718],seed[2983],seed[2685],seed[1730],seed[3028],seed[3784],seed[1376],seed[1414],seed[1770],seed[2648],seed[1572],seed[597],seed[3740],seed[2298],seed[3673],seed[3603],seed[2521],seed[3843],seed[3407],seed[1759],seed[46],seed[2751],seed[2147],seed[1897],seed[2978],seed[3437],seed[448],seed[2153],seed[2100],seed[1160],seed[1382],seed[2614],seed[3251],seed[3277],seed[3990],seed[3135],seed[601],seed[1251],seed[617],seed[789],seed[1211],seed[4050],seed[716],seed[2296],seed[2184],seed[3347],seed[2288],seed[3889],seed[4064],seed[730],seed[207],seed[486],seed[1564],seed[555],seed[1407],seed[155],seed[1976],seed[682],seed[2675],seed[1655],seed[3621],seed[1206],seed[491],seed[3453],seed[3789],seed[1005],seed[3528],seed[2750],seed[261],seed[1043],seed[3232],seed[1970],seed[3947],seed[2370],seed[2941],seed[333],seed[1519],seed[1510],seed[3156],seed[2563],seed[1848],seed[1269],seed[947],seed[3907],seed[902],seed[3931],seed[509],seed[2929],seed[778],seed[1296],seed[1701],seed[2901],seed[982],seed[3202],seed[2152],seed[1902],seed[198],seed[2062],seed[2844],seed[2140],seed[3520],seed[3688],seed[784],seed[2308],seed[3053],seed[382],seed[1431],seed[2723],seed[1529],seed[1997],seed[3479],seed[183],seed[2619],seed[3509],seed[723],seed[1645],seed[1007],seed[1194],seed[1168],seed[2086],seed[308],seed[1889],seed[341],seed[2222],seed[2213],seed[1430],seed[780],seed[1666],seed[3412],seed[3067],seed[1209],seed[3766],seed[662],seed[3385],seed[1958],seed[492],seed[695],seed[1561],seed[1397],seed[1371],seed[1754],seed[108],seed[424],seed[604],seed[2762],seed[2402],seed[3712],seed[3138],seed[1637],seed[175],seed[900],seed[4004],seed[2584],seed[2314],seed[1062],seed[1399],seed[293],seed[2914],seed[2161],seed[3886],seed[980],seed[3370],seed[4065],seed[1245],seed[158],seed[521],seed[130],seed[2212],seed[1110],seed[3307],seed[3682],seed[3660],seed[2855],seed[254],seed[2609],seed[9],seed[2937],seed[3454],seed[2861],seed[3636],seed[758],seed[511],seed[3519],seed[527],seed[422],seed[1339],seed[573],seed[2395],seed[299],seed[2165],seed[3853],seed[3567],seed[3937],seed[1347],seed[3661],seed[389],seed[3267],seed[2096],seed[1815],seed[1498],seed[2650],seed[794],seed[3387],seed[3271],seed[3882],seed[1813],seed[2627],seed[2657],seed[3086],seed[2838],seed[2730],seed[2210],seed[3494],seed[1299],seed[1357],seed[202],seed[322],seed[420],seed[2134],seed[2012],seed[3273],seed[1349],seed[2965],seed[51],seed[2935],seed[74],seed[967],seed[1212],seed[3457],seed[2172],seed[1023],seed[1745],seed[2342],seed[1996],seed[2879],seed[3901],seed[2185],seed[154],seed[85],seed[3078],seed[2214],seed[215],seed[3570],seed[2728],seed[1530],seed[2175],seed[1122],seed[3809],seed[1396],seed[3476],seed[2257],seed[3652],seed[1622],seed[848],seed[1180],seed[3339],seed[1022],seed[2275],seed[3912],seed[1141],seed[2158],seed[2238],seed[289],seed[2355],seed[569],seed[3217],seed[3506],seed[1649],seed[565],seed[2871],seed[1142],seed[1845],seed[2490],seed[2235],seed[1364],seed[1668],seed[2125],seed[2323],seed[3213],seed[1085],seed[3617],seed[318],seed[994],seed[230],seed[3909],seed[2516],seed[2114],seed[415],seed[632],seed[909],seed[951],seed[1317],seed[1964],seed[2203],seed[649],seed[645],seed[1948],seed[1176],seed[3706],seed[1583],seed[1352],seed[3609],seed[1960],seed[3753],seed[1609],seed[2806],seed[3128],seed[460],seed[4042],seed[3736],seed[953],seed[2899],seed[3869],seed[2121],seed[219],seed[1385],seed[3994],seed[103],seed[1837],seed[88],seed[885],seed[3503],seed[2766],seed[3633],seed[4071],seed[410],seed[2888],seed[2961],seed[157],seed[567],seed[2290],seed[523],seed[3285],seed[641],seed[457],seed[160],seed[400],seed[223],seed[2434],seed[1586],seed[3689],seed[1779],seed[3101],seed[4017],seed[3493],seed[1593],seed[3950],seed[2705],seed[136],seed[2108],seed[2351],seed[786],seed[2072],seed[2956],seed[924],seed[3906],seed[2958],seed[1823],seed[2880],seed[2683],seed[1767],seed[2854],seed[3112],seed[2039],seed[1500],seed[2835],seed[271],seed[2091],seed[1766],seed[2664],seed[561],seed[2805],seed[3207],seed[530],seed[3619],seed[1624],seed[2302],seed[1097],seed[1629],seed[248],seed[19],seed[2892],seed[2803],seed[2549],seed[2135],seed[1053],seed[1320],seed[3548],seed[1291],seed[628],seed[1157],seed[3697],seed[2483],seed[1466],seed[2939],seed[3296],seed[1208],seed[816],seed[547],seed[1654],seed[177],seed[918],seed[2923],seed[2389],seed[996],seed[485],seed[732],seed[2727],seed[1746],seed[4095],seed[3471],seed[3835],seed[972],seed[3829],seed[1824],seed[529],seed[2863],seed[2515],seed[1453],seed[73],seed[394],seed[4053],seed[1771],seed[3513],seed[4015],seed[3206],seed[390],seed[1205],seed[3191],seed[3516],seed[253],seed[737],seed[3921],seed[2885],seed[1204],seed[2128],seed[2057],seed[2647],seed[2503],seed[3171],seed[3709],seed[2967],seed[2597],seed[3733],seed[1031],seed[680],seed[1484],seed[164],seed[2010],seed[3504],seed[3033],seed[2702],seed[3464],seed[440],seed[206],seed[971],seed[830],seed[575],seed[292],seed[2847],seed[1018],seed[993],seed[912],seed[592],seed[3338],seed[1661],seed[4067],seed[3978],seed[1667],seed[2966],seed[316],seed[3137],seed[3648],seed[4036],seed[89],seed[3314],seed[2478],seed[3642],seed[3678],seed[1086],seed[2712],seed[2295],seed[3438],seed[2862],seed[3954],seed[1330],seed[3258],seed[2240],seed[2348],seed[872],seed[1715],seed[1246],seed[2102],seed[1546],seed[3113],seed[1720],seed[52],seed[1452],seed[4052],seed[775],seed[2662],seed[3898],seed[1064],seed[210],seed[489],seed[1136],seed[2560],seed[3325],seed[1116],seed[311],seed[3490],seed[2004],seed[2332],seed[965],seed[2263],seed[3189],seed[2535],seed[1181],seed[2189],seed[1354],seed[3379],seed[2453],seed[3220],seed[2799],seed[2786],seed[1615],seed[2668],seed[2477],seed[1446],seed[487],seed[2949],seed[1955],seed[1461],seed[3797],seed[233],seed[2069],seed[2920],seed[2306],seed[1680],seed[2607],seed[3293],seed[2473],seed[2637],seed[2573],seed[3359],seed[3115],seed[3641],seed[570],seed[3272],seed[456],seed[2347],seed[709],seed[1153],seed[2593],seed[1838],seed[399],seed[3276],seed[2699],seed[1036],seed[3803],seed[2928],seed[8],seed[1381],seed[1095],seed[3545],seed[3175],seed[1513],seed[442],seed[3943],seed[2718],seed[3139],seed[2532],seed[3160],seed[781],seed[1081],seed[823],seed[2669],seed[958],seed[3009],seed[788],seed[3948],seed[1696],seed[2460],seed[1221],seed[1263],seed[704],seed[3914],seed[1731],seed[117],seed[3341],seed[1282],seed[3110],seed[1140],seed[3505],seed[228],seed[4058],seed[1589],seed[679],seed[1869],seed[1576],seed[2737],seed[2865],seed[2527],seed[3436],seed[423],seed[2789],seed[3245],seed[538],seed[3125],seed[3243],seed[1236],seed[519],seed[3036],seed[2747],seed[3897],seed[1984],seed[710],seed[1285],seed[3211],seed[2782],seed[2426],seed[2580],seed[1014],seed[4045],seed[1459],seed[837],seed[124],seed[1679],seed[331],seed[3116],seed[1550],seed[822],seed[1538],seed[2623],seed[2058],seed[3507],seed[344],seed[3363],seed[1855],seed[25],seed[3888],seed[3153],seed[3380],seed[3925],seed[4007],seed[1517],seed[3345],seed[1785],seed[542],seed[417],seed[3604],seed[3157],seed[76],seed[3499],seed[1863],seed[13],seed[633],seed[1473],seed[2542],seed[67],seed[1728],seed[1856],seed[2216],seed[3404],seed[329],seed[1947],seed[2595],seed[335],seed[1794],seed[2231],seed[1692],seed[1093],seed[2280],seed[1108],seed[1173],seed[1651],seed[1326],seed[1297],seed[771],seed[3971],seed[143],seed[883],seed[3854],seed[2823],seed[1698],seed[1019],seed[2821],seed[502],seed[3615],seed[2377],seed[2282],seed[4000],seed[3440],seed[476],seed[2368],seed[3095],seed[2007],seed[1543],seed[243],seed[3722],seed[2895],seed[403],seed[3281],seed[1893],seed[3366],seed[3981],seed[3832],seed[225],seed[4023],seed[3495],seed[2707],seed[847],seed[2617],seed[3234],seed[60],seed[2971],seed[990],seed[1230],seed[2437],seed[2363],seed[3039],seed[4076],seed[4019],seed[113],seed[747],seed[2759],seed[640],seed[1542],seed[3424],seed[1226],seed[941],seed[3614],seed[3685],seed[1750],seed[893],seed[3342],seed[1697],seed[2973],seed[2379],seed[2466],seed[4027],seed[2499],seed[239],seed[104],seed[2903],seed[234],seed[2482],seed[1045],seed[1791],seed[1432],seed[1709],seed[3561],seed[1532],seed[700],seed[2463],seed[2725],seed[4094],seed[365],seed[2136],seed[2447],seed[285],seed[2469],seed[669],seed[2876],seed[1826],seed[745],seed[3330],seed[862],seed[378],seed[1096],seed[1986],seed[1469],seed[1336],seed[3391],seed[678],seed[4006],seed[2180],seed[3131],seed[200],seed[2415],seed[1101],seed[452],seed[1126],seed[841],seed[2846],seed[1415],seed[696],seed[1207],seed[2760],seed[2160],seed[310],seed[4056],seed[1999],seed[798],seed[1858],seed[357],seed[3526],seed[1665],seed[1919],seed[634],seed[3515],seed[2663],seed[3237],seed[648],seed[2975],seed[1272],seed[3775],seed[224],seed[2250],seed[1507],seed[4003],seed[1425],seed[3899],seed[1951],seed[3840],seed[2051],seed[2101],seed[3389],seed[2801],seed[3275],seed[1935],seed[2429],seed[549],seed[2922],seed[1198],seed[2038],seed[2026],seed[1197],seed[4010],seed[82],seed[690],seed[77],seed[435],seed[2470],seed[3579],seed[1408],seed[2673],seed[3744],seed[1429],seed[2770],seed[3127],seed[2398],seed[677],seed[2646],seed[1151],seed[3824],seed[36],seed[4079],seed[1312],seed[2601],seed[2391],seed[624],seed[336],seed[2656],seed[3554],seed[1660],seed[2860],seed[106],seed[3560],seed[708],seed[2566],seed[2757],seed[3798],seed[120],seed[3238],seed[2365],seed[3502],seed[3032],seed[2050],seed[3332],seed[3195],seed[2107],seed[2392],seed[2090],seed[23],seed[184],seed[3406],seed[1894],seed[1805],seed[3932],seed[3764],seed[2710],seed[1836],seed[2232],seed[275],seed[3668],seed[2740],seed[1941],seed[3591],seed[861],seed[540],seed[231],seed[3517],seed[4082],seed[2186],seed[1975],seed[3483],seed[3107],seed[1934],seed[916],seed[1844],seed[201],seed[2319],seed[3382],seed[884],seed[3320],seed[3872],seed[105],seed[2817],seed[3836],seed[2583],seed[2412],seed[1772],seed[831],seed[141],seed[3821],seed[1670],seed[3018],seed[2143],seed[1891],seed[2028],seed[1069],seed[3123],seed[2955],seed[1909],seed[3247],seed[2701],seed[2046],seed[4016],seed[2825],seed[1169],seed[1188],seed[3655],seed[797],seed[2179],seed[2061],seed[2413],seed[3555],seed[3208],seed[220],seed[3696],seed[929],seed[4048],seed[688],seed[251],seed[2097],seed[4033],seed[1384],seed[1795],seed[2495],seed[1174],seed[3260],seed[1928],seed[3420],seed[1783],seed[65],seed[2795],seed[2665],seed[3224],seed[2094],seed[1088],seed[528],seed[1398],seed[3169],seed[2582],seed[1601],seed[3558],seed[3178],seed[1927],seed[1711],seed[1274],seed[843],seed[3346],seed[1041],seed[579],seed[804],seed[2635],seed[1907],seed[2845],seed[653],seed[3527],seed[2224],seed[3003],seed[599],seed[466],seed[937],seed[3769],seed[1026],seed[2278],seed[1872],seed[2947],seed[3394],seed[1133],seed[2171],seed[431],seed[2170],seed[3933],seed[3060],seed[1575],seed[583],seed[375],seed[404],seed[3691],seed[956],seed[2887],seed[2373],seed[407],seed[3073],seed[2514],seed[332],seed[3934],seed[49],seed[266],seed[2011],seed[3825],seed[821],seed[1784],seed[3540],seed[718],seed[2401],seed[2792],seed[342],seed[1659],seed[1039],seed[1954],seed[369],seed[3396],seed[3158],seed[3108],seed[1977],seed[12],seed[3757],seed[891],seed[3235],seed[805],seed[2918],seed[1061],seed[2643],seed[672],seed[811],seed[3362],seed[1420],seed[286],seed[212],seed[2993],seed[1258],seed[955],seed[465],seed[3525],seed[2713],seed[844],seed[3857],seed[1071],seed[1146],seed[1387],seed[2076],seed[2872],seed[808],seed[1877],seed[3827],seed[2571],seed[3063],seed[392],seed[2547],seed[4088],seed[2997],seed[2802],seed[196],seed[1663],seed[3057],seed[3430],seed[3720],seed[40],seed[3632],seed[3628],seed[1228],seed[2852],seed[3000],seed[666],seed[1224],seed[1641],seed[2704],seed[3596],seed[515],seed[3304],seed[2192],seed[2071],seed[2324],seed[2018],seed[3481],seed[3855],seed[413],seed[2940],seed[2843],seed[4032],seed[1604],seed[2790],seed[55],seed[1918],seed[1454],seed[2708],seed[3222],seed[3278],seed[548],seed[1683],seed[371],seed[4063],seed[1],seed[1677],seed[1717],seed[2080],seed[3608],seed[2896],seed[2145],seed[2444],seed[3368],seed[2118],seed[623],seed[3957],seed[1778],seed[1074],seed[3223],seed[3069],seed[3936],seed[921],seed[21],seed[1293],seed[2113],seed[3928],seed[2518],seed[2869],seed[3643],seed[1082],seed[2042],seed[881],seed[2558],seed[482],seed[2574],seed[1578],seed[2645],seed[1551],seed[1648],seed[724],seed[139],seed[3480],seed[2191],seed[3445],seed[533],seed[2731],seed[3257],seed[612],seed[1994],seed[2139],seed[731],seed[3002],seed[2253],seed[2181],seed[2743],seed[796],seed[550],seed[3197],seed[740],seed[1913],seed[2546],seed[1276],seed[2837],seed[987],seed[536],seed[759],seed[1424],seed[144],seed[770],seed[169],seed[2268],seed[453],seed[2411],seed[2251],seed[3622],seed[43],seed[2606],seed[932],seed[2047],seed[3261],seed[1761],seed[588],seed[1985],seed[580],seed[2906],seed[3219],seed[2227],seed[1887],seed[2052],seed[2716],seed[1137],seed[2099],seed[2427],seed[3626],seed[4008],seed[1528],seed[2040],seed[3795],seed[908],seed[1524],seed[1266],seed[2089],seed[3162],seed[2828],seed[806],seed[2449],seed[2926],seed[1652],seed[112],seed[2375],seed[1865],seed[3814],seed[2894],seed[674],seed[2310],seed[1159],seed[2327],seed[2996],seed[3765],seed[735],seed[3724],seed[1467],seed[1416],seed[2953],seed[3731],seed[1154],seed[3637],seed[2221],seed[3917],seed[743],seed[2959],seed[2649],seed[1494],seed[3601],seed[3180],seed[2423],seed[2334],seed[767],seed[2618],seed[850],seed[1201],seed[1118],seed[3521],seed[1373],seed[2273],seed[3274],seed[1705],seed[1850],seed[564],seed[2689],seed[3910],seed[3828],seed[1802],seed[3951],seed[115],seed[147],seed[1769],seed[3375],seed[3598],seed[4005],seed[3692],seed[1688],seed[2019],seed[1816],seed[2318],seed[3093],seed[114],seed[1318],seed[3704],seed[2505],seed[3042],seed[3799],seed[1890],seed[3998],seed[1541],seed[3987],seed[2900],seed[2380],seed[2672],seed[2151],seed[2839],seed[3826],seed[1922],seed[3877],seed[127],seed[1789],seed[1614],seed[3164],seed[2556],seed[2927],seed[657],seed[2367],seed[81],seed[3543],seed[3941],seed[3145],seed[324],seed[4068],seed[1669],seed[3589],seed[501],seed[2305],seed[1215],seed[2182],seed[2098],seed[178],seed[2496],seed[2487],seed[4092],seed[2024],seed[2698],seed[1516],seed[2283],seed[2265],seed[2753],seed[2336],seed[1574],seed[2311],seed[545],seed[4046],seed[1451],seed[2462],seed[1884],seed[2857],seed[3707],seed[1846],seed[3865],seed[3462],seed[170],seed[1747],seed[3126],seed[1582],seed[1762],seed[673],seed[952],seed[1441],seed[111],seed[3737],seed[80],seed[2919],seed[2127],seed[2576],seed[6],seed[1072],seed[1010],seed[3913],seed[946],seed[2043],seed[2729],seed[277],seed[2122],seed[1867],seed[3742],seed[205],seed[84],seed[3225],seed[685],seed[1639],seed[3097],seed[2765],seed[1162],seed[216],seed[865],seed[358],seed[1623],seed[2141],seed[915],seed[2027],seed[877],seed[4039],seed[276],seed[2798],seed[1694],seed[295],seed[1506],seed[3204],seed[93],seed[2312],seed[2079],seed[2016],seed[2776],seed[398],seed[3360],seed[4072],seed[1793],seed[3241],seed[1636],seed[3012],seed[2432],seed[3734],seed[1981],seed[3647],seed[31],seed[1428],seed[832],seed[3199],seed[1926],seed[3443],seed[2316],seed[2533],seed[3315],seed[3151],seed[637],seed[3927],seed[734],seed[3068],seed[3659],seed[1040],seed[3967],seed[2344],seed[868],seed[1368],seed[3161],seed[1184],seed[896],seed[1650],seed[2651],seed[1565],seed[554],seed[833],seed[2162],seed[562],seed[572],seed[2048],seed[1768],seed[2671],seed[1389],seed[2946],seed[2281],seed[1075],seed[522],seed[1275],seed[3284],seed[1308],seed[1833],seed[1931],seed[1148],seed[2575],seed[3433],seed[3122],seed[907],seed[684],seed[541],seed[3300],seed[3035],seed[1254],seed[736],seed[2824],seed[1818],seed[2562],seed[374],seed[2301],seed[2372],seed[2758],seed[2544],seed[4020],seed[2362],seed[574],seed[3231],seed[2764],seed[3085],seed[1870],seed[875],seed[764],seed[1904],seed[1673],seed[566],seed[1400],seed[3719],seed[871],seed[2613],seed[1883],seed[1278],seed[193],seed[2693],seed[2243],seed[1952],seed[991],seed[2523],seed[4024],seed[2554],seed[2615],seed[1448],seed[2218],seed[934],seed[3045],seed[3102],seed[2706],seed[2060],seed[1812],seed[1046],seed[3552],seed[3333],seed[4025],seed[1147],seed[1625],seed[2994],seed[935],seed[2884],seed[1968],seed[2735],seed[857],seed[4040],seed[2970],seed[512],seed[3830],seed[1643],seed[2220],seed[211],seed[763],seed[3254],seed[2260],seed[2811],seed[2315],seed[3316],seed[984],seed[1238],seed[1163],seed[161],seed[2632],seed[2359],seed[1232],seed[1322],seed[107],seed[3027],seed[3542],seed[867],seed[499],seed[4051],seed[1503],seed[1288],seed[3962],seed[1050],seed[1035],seed[3323],seed[444],seed[1713],seed[2188],seed[3472],seed[2721],seed[1886],seed[1658],seed[3061],seed[1504],seed[596],seed[3079],seed[1840],seed[1161],seed[3313],seed[1068],seed[1348],seed[3966],seed[819],seed[1949],seed[4014],seed[1488],seed[1882],seed[1143],seed[3915],seed[2123],seed[1367],seed[2781],seed[370],seed[1776],seed[1827],seed[1773],seed[3781],seed[2769],seed[2777],seed[98],seed[2506],seed[2406],seed[2744],seed[1920],seed[1515],seed[438],seed[1612],seed[3823],seed[1721],seed[1025],seed[2196],seed[1411],seed[729],seed[3295],seed[3804],seed[2755],seed[3758],seed[345],seed[1092],seed[2115],seed[38],seed[3788],seed[2780],seed[615],seed[376],seed[2335],seed[2405],seed[1595],seed[2441],seed[1422],seed[1874],seed[2536],seed[1950],seed[3187],seed[1522],seed[3701],seed[4002],seed[2297],seed[1803],seed[320],seed[1687],seed[4080],seed[167],seed[361],seed[2567],seed[2629],seed[3328],seed[87],seed[3754],seed[518],seed[1403],seed[897],seed[50],seed[469],seed[2692],seed[1881],seed[3062],seed[1724],seed[1063],seed[3147],seed[3666],seed[1421],seed[504],seed[472],seed[3538],seed[505],seed[1483],seed[2891],seed[284],seed[4029],seed[195],seed[2974],seed[3263],seed[4077],seed[1440],seed[3968],seed[762],seed[2577],seed[2608],seed[3422],seed[2797],seed[57],seed[3856],seed[53],seed[3104],seed[756],seed[468],seed[2654],seed[2522],seed[1868],seed[3469],seed[279],seed[1223],seed[3894],seed[3774],seed[278],seed[1733],seed[459],seed[560],seed[379],seed[303],seed[2480],seed[2049],seed[3386],seed[2526],seed[3801],seed[3324],seed[3419],seed[1509],seed[2564],seed[1710],seed[631],seed[2386],seed[3813],seed[3559],seed[1257],seed[3565],seed[981],seed[1457],seed[817],seed[1301],seed[1132],seed[2002],seed[3343],seed[3159],seed[1995],seed[3488],seed[859],seed[2326],seed[1618],seed[1906],seed[1359],seed[1073],seed[1443],seed[373],seed[3911],seed[3983],seed[3473],seed[1495],seed[3999],seed[2006],seed[719],seed[3859],seed[325],seed[686],seed[1716],seed[2980],seed[714],seed[1084],seed[3264],seed[3352],seed[3920],seed[425],seed[235],seed[3748],seed[3716],seed[3004],seed[3305],seed[1600],seed[1485],seed[1241],seed[1978],seed[354],seed[559],seed[1972],seed[3050],seed[280],seed[1946],seed[3568],seed[751],seed[3790],seed[1012],seed[1988],seed[1860],seed[887],seed[2309],seed[349],seed[1944],seed[481],seed[3331],seed[3183],seed[1127],seed[3327],seed[1051],seed[3358],seed[1765],seed[1222],seed[2303],seed[1956],seed[2788],seed[1294],seed[3811],seed[728],seed[713],seed[2734],seed[939],seed[2594],seed[445],seed[705],seed[2603],seed[3762],seed[1192],seed[498],seed[3923],seed[910],seed[944],seed[10],seed[2599],seed[471],seed[1214],seed[1052],seed[2321],seed[3065],seed[977],seed[2631],seed[989],seed[1243],seed[2410],seed[2378],seed[3550],seed[2904],seed[2293],seed[1939],seed[2794],seed[1774],seed[1409],seed[281],seed[45],seed[1809],seed[2440],seed[663],seed[3532],seed[26],seed[1410],seed[894],seed[2957],seed[1478],seed[246],seed[1463],seed[2659],seed[3945],seed[1932],seed[1702],seed[2394],seed[2031],seed[904],seed[2357],seed[2077],seed[517],seed[1402],seed[3092],seed[3600],seed[3592],seed[241],seed[1374],seed[3392],seed[1689],seed[2497],seed[2197],seed[125],seed[3980],seed[2459],seed[405],seed[1959],seed[3868],seed[3006],seed[1417],seed[1632],seed[3761],seed[2381],seed[119],seed[1905],seed[388],seed[1549],seed[122],seed[1908],seed[309],seed[2337],seed[3049],seed[1725],seed[2512],seed[3020],seed[785],seed[406],seed[610],seed[537],seed[2464],seed[3306],seed[750],seed[2126],seed[2073],seed[2258],seed[3749],seed[2889],seed[3776],seed[699],seed[2754],seed[886],seed[1130],seed[2703],seed[301],seed[56],seed[174],seed[2856],seed[37],seed[2655],seed[1255],seed[1165],seed[1302],seed[2924],seed[17],seed[2746],seed[1379],seed[1900],seed[172],seed[1866],seed[434],seed[2552],seed[2485],seed[942],seed[3582],seed[1796],seed[644],seed[2284],seed[1547],seed[973],seed[2361],seed[914],seed[742],seed[131],seed[1569],seed[3099],seed[3955],seed[1178],seed[2105],seed[2510],seed[3432],seed[621],seed[2963],seed[854],seed[1518],seed[3090],seed[3756],seed[2084],seed[2032],seed[2778],seed[232],seed[3470],seed[2622],seed[1247],seed[1129],seed[3985],seed[446],seed[3970],seed[2684],seed[820],seed[3074],seed[2779],seed[3026],seed[834],seed[2408],seed[3881],seed[2358],seed[2146],seed[1033],seed[1098],seed[24],seed[1358],seed[1365],seed[576],seed[3862],seed[2059],seed[2202],seed[2030],seed[264],seed[3739],seed[2286],seed[1631],seed[2467],seed[2819],seed[3408],seed[1591],seed[2866],seed[3782],seed[2717],seed[2356],seed[2667],seed[3512],seed[658],seed[1471],seed[3892],seed[1388],seed[1008],seed[3083],seed[4001],seed[1321],seed[3322],seed[1057],seed[1311],seed[3082],seed[3908],seed[441],seed[3043],seed[1590],seed[3040],seed[2620],seed[3864],seed[3848],seed[477],seed[1880],seed[2353],seed[1987],seed[3665],seed[930],seed[1544],seed[1465],seed[3721],seed[664],seed[247],seed[3037],seed[3845],seed[110],seed[1315],seed[3188],seed[4090],seed[83],seed[128],seed[3723],seed[860],seed[3553],seed[66],seed[557],seed[838],seed[563],seed[3109],seed[1164],seed[2498],seed[3566],seed[3335],seed[3141],seed[1851],seed[1775],seed[409],seed[3198],seed[1914],seed[2219],seed[99],seed[1248],seed[488],seed[1751],seed[1316],seed[3373],seed[532],seed[287],seed[578],seed[1496],seed[3610],seed[2148],seed[1034],seed[265],seed[3866],seed[754],seed[898],seed[2587],seed[2149],seed[3735],seed[2513],seed[3024],seed[2796],seed[1447],seed[29],seed[1286],seed[2461],seed[1917],seed[3885],seed[1427],seed[1657],seed[3533],seed[1021],seed[1264],seed[3240],seed[2199],seed[3991],seed[1455],seed[1579],seed[451],seed[2504],seed[20],seed[2768],seed[1611],seed[156],seed[2132],seed[3265],seed[3226],seed[2832],seed[3303],seed[1307],seed[3310],seed[1991],seed[3193],seed[3094],seed[1267],seed[3140],seed[1329],seed[3564],seed[3114],seed[2117],seed[3562],seed[2183],seed[873],seed[1965],seed[1607],seed[2785],seed[259],seed[2065],seed[799],seed[2244],seed[1167],seed[62],seed[1690],seed[3919],seed[1971],seed[3658],seed[2984],seed[948],seed[765],seed[3354],seed[2726],seed[643],seed[2041],seed[1501],seed[2990],seed[1259],seed[3677],seed[2831],seed[191],seed[4091],seed[1090],seed[1545],seed[760],seed[701],seed[2211],seed[4086],seed[42],seed[2813],seed[2596],seed[2666],seed[3942],seed[1011],seed[825],seed[923],seed[2938],seed[3871],seed[2660],seed[1378],seed[462],seed[3551],seed[1933],seed[3249],seed[1249],seed[4041],seed[801],seed[779],seed[4078],seed[47],seed[2881],seed[1295],seed[3606],seed[1135],seed[3046],seed[3100],seed[199],seed[826],seed[1854],seed[2157],seed[2822],seed[1674],seed[294],seed[3172],seed[1548],seed[3047],seed[2875],seed[2078],seed[2589],seed[3819],seed[1628],seed[2442],seed[3715],seed[2068],seed[1076],seed[2652],seed[386],seed[2960],seed[3587],seed[63],seed[2772],seed[41],seed[2676],seed[450],seed[1490],seed[109],seed[306],seed[2252],seed[691],seed[3405],seed[366],seed[534],seed[1145],seed[3662],seed[3398],seed[1969],seed[2551],seed[1675],seed[1508],seed[2245],seed[1213],seed[256],seed[1094],seed[608],seed[3858],seed[3279],seed[368],seed[2989],seed[3717],seed[1512],seed[1562],seed[3725],seed[2952],seed[1152],seed[2045],seed[815],seed[2349],seed[2167],seed[938],seed[3337],seed[3447],seed[3729],seed[960],seed[302],seed[190],seed[2827],seed[1584],seed[1640],seed[702],seed[203],seed[726],seed[2354],seed[3732],seed[793],seed[2396],seed[3524],seed[879],seed[795],seed[2886],seed[2109],seed[3444],seed[3572],seed[851],seed[707],seed[48],seed[3602],seed[229],seed[3318],seed[3613],seed[2277],seed[2592],seed[2259],seed[1003],seed[3428],seed[3989],seed[2131],seed[1819],seed[347],seed[2083],seed[3841],seed[2023],seed[1361],seed[2830],seed[571],seed[3687],seed[2092],seed[911],seed[221],seed[1536],seed[3575],seed[463],seed[3403],seed[2330],seed[3150],seed[1790],seed[1350],seed[496],seed[2],seed[3072],seed[4028],seed[722],seed[455],seed[1139],seed[1177],seed[3771],seed[3796],seed[3863],seed[1131],seed[2384],seed[2686],seed[2748],seed[217],seed[1760],seed[1059],seed[2409],seed[1029],seed[1753],seed[2093],seed[1990],seed[3088],seed[1338],seed[890],seed[2393],seed[3805],seed[2067],seed[314],seed[3259],seed[556],seed[3926],seed[3620],seed[3767],seed[2194],seed[1191],seed[1945],seed[3077],seed[3590],seed[568],seed[1525],seed[3946],seed[1170],seed[433],seed[142],seed[3630],seed[1438],seed[3569],seed[2176],seed[1231],seed[4055],seed[1610],seed[3807],seed[2407],seed[2472],seed[1567],seed[3786],seed[1656],seed[524],seed[551],seed[15],seed[3397],seed[1458],seed[1817],seed[408],seed[151],seed[414],seed[3329],seed[2075],seed[263],seed[2417],seed[2269],seed[3938],seed[3728],seed[2085],seed[3873],seed[3054],seed[393],seed[584],seed[3842],seed[2925],seed[3144],seed[1185],seed[3194],seed[3675],seed[2809],seed[28],seed[3297],seed[2168],seed[1718],seed[1493],seed[255],seed[995],seed[2908],seed[602],seed[2360],seed[1048],seed[2020],seed[2029],seed[2742],seed[3791],seed[2968],seed[4022],seed[979],seed[2207],seed[639],seed[1309],seed[1186],seed[1091],seed[2366],seed[1107],seed[118],seed[1028],seed[1621],seed[1001],seed[3402],seed[2022],seed[3173],seed[1744],seed[149],seed[2420],seed[1531],seed[159],seed[3168],seed[4069],seed[1182],seed[2229],seed[1682],seed[2400],seed[2475],seed[2155],seed[1892],seed[1303],seed[2364],seed[137],seed[2907],seed[2350],seed[3401],seed[1712],seed[508],seed[3434],seed[2003],seed[102],seed[359],seed[1000],seed[1190],seed[4013],seed[3288],seed[1752],seed[3940],seed[3657],seed[2451],seed[2541],seed[2833],seed[866],seed[2661],seed[1380],seed[3850],seed[1520],seed[4047],seed[478],seed[2545],seed[2088],seed[1616],seed[943],seed[842],seed[1613],seed[968],seed[2962],seed[3986],seed[2341],seed[1366],seed[3686],seed[283],seed[5],seed[2557],seed[2910],seed[1873],seed[3482],seed[3356],seed[1916],seed[3361],seed[2005],seed[2853],seed[227],seed[1810],seed[1570],seed[2205],seed[3124],seed[3959],seed[1273],seed[3884],seed[3051],seed[2715],seed[3022],seed[2195],seed[2142],seed[525],seed[3847],seed[3376],seed[470],seed[976],seed[1808],seed[3583],seed[2431],seed[2130],seed[1553],seed[2502],seed[411],seed[2678],seed[635],seed[603],seed[1814],seed[1878],seed[3627],seed[2274],seed[2438],seed[3477],seed[1435],seed[3531],seed[1327],seed[2773],seed[64],seed[3253],seed[2333],seed[1699],seed[3233],seed[3336],seed[741],seed[1849],seed[3816],seed[1523],seed[2285],seed[3446],seed[1439],seed[58],seed[1749],seed[3417],seed[1842],seed[3547],seed[3918],seed[3181],seed[1957],seed[1256],seed[484],seed[2385],seed[3759],seed[3388],seed[1179],seed[2818],seed[4021],seed[1862],seed[3586],seed[2816],seed[3423],seed[3084],seed[240],seed[1449],seed[3780],seed[213],seed[3646],seed[493],seed[2931],seed[3034],seed[464],seed[1821],seed[2267],seed[86],seed[630],seed[3400],seed[2540],seed[1331],seed[3413],seed[298],seed[296],seed[2680],seed[945],seed[3890],seed[864],seed[1277],seed[267],seed[3746],seed[3680],seed[1961],seed[2930],seed[2912],seed[2793],seed[1089],seed[3087],seed[2340],seed[2403],seed[2812],seed[2013],seed[126],seed[3979],seed[1300],seed[1346],seed[1150],seed[2255],seed[1585],seed[1187],seed[3653],seed[1464],seed[1634],seed[1037],seed[2642],seed[1505],seed[899],seed[2479],seed[1499],seed[3963],seed[2111],seed[3793],seed[339],seed[1895],seed[1183],seed[882],seed[3229],seed[1103],seed[3317],seed[2991],seed[2578],seed[1620],seed[3439],seed[1401],seed[3997],seed[2842],seed[4087],seed[3710],seed[16],seed[30],seed[3255],seed[922],seed[2489],seed[237],seed[790],seed[3891],seed[4026],seed[3299],seed[1289],seed[2374],seed[439],seed[2008],seed[852],seed[1676],seed[1383],seed[2581],seed[395],seed[1535],seed[2864],seed[4059],seed[304],seed[132],seed[1460],seed[3992],seed[313],seed[1831],seed[1587],seed[3849],seed[100],seed[4081],seed[687],seed[2492],seed[1811],seed[3511],seed[1369],seed[3014],seed[1723],seed[949],seed[2591],seed[3117],seed[44],seed[2995],seed[176],seed[1437],seed[1912],seed[2543],seed[2064],seed[419],seed[454],seed[3492],seed[1708],seed[1521],seed[1847],seed[3574],seed[2439],seed[1047],seed[3611],seed[3236],seed[2714],seed[2137],seed[2500],seed[1386],seed[428],seed[2081],seed[2346],seed[2763],seed[249],seed[260],seed[1729],seed[2369],seed[269],seed[3218],seed[582],seed[2644],seed[757],seed[3977],seed[2588],seed[2877],seed[2234],seed[3964],seed[1334],seed[1283],seed[905],seed[1915],seed[2242],seed[3817],seed[2455],seed[2736],seed[1233],seed[2936],seed[2690],seed[2488],seed[581],seed[3778],seed[1896],seed[1351],seed[348],seed[3016],seed[1859],seed[1227],seed[783],seed[3179],seed[810],seed[2272],seed[3844],seed[1020],seed[2430],seed[591],seed[613],seed[1822],seed[4093],seed[1344],seed[4044],seed[2352],seed[2021],seed[2074],seed[1189],seed[2909],seed[2294],seed[3038],seed[1577],seed[2579],seed[1111],seed[3001],seed[1042],seed[619],seed[3132],seed[650],seed[2169],seed[3041],seed[1099],seed[2201],seed[2313],seed[2494],seed[78],seed[3537],seed[2230],seed[3763],seed[818],seed[2981],seed[3585],seed[926],seed[4037],seed[97],seed[660],seed[92],seed[855],seed[401],seed[3895],seed[2870],seed[1973],seed[3852],seed[903],seed[928],seed[1080],seed[1596],seed[917],seed[2390],seed[1588],seed[3378],seed[1839],seed[494],seed[2299],seed[2628],seed[3426],seed[3390],seed[611],seed[836],seed[2977],seed[739],seed[3549],seed[2150],seed[2840],seed[1426],seed[2979],seed[2082],seed[1196],seed[3010],seed[3015],seed[3308],seed[1125],seed[3081],seed[2720],seed[2911],seed[2036],seed[3594],seed[2807],seed[2988],seed[787],seed[2215],seed[396],seed[1533],seed[3381],seed[1719],seed[2550],seed[1149],seed[2943],seed[1804],seed[372],seed[2964],seed[2921],seed[4038],seed[3523],seed[473],seed[27],seed[1756],seed[3121],seed[1335],seed[1216],seed[3563],seed[166],seed[288],seed[2711],seed[3867],seed[1172],seed[1857],seed[307],seed[2416],seed[2397],seed[2572],seed[3802],seed[402],seed[1864],seed[1260],seed[242],seed[2733],seed[3466],seed[479],seed[768],seed[3738],seed[2836],seed[1055],seed[1633],seed[2343],seed[2537],seed[3768],seed[3212],seed[2917],seed[627],seed[2610],seed[3205],seed[188],seed[2586],seed[920],seed[1560],seed[3752],seed[870],seed[1328],seed[1899],seed[1843],seed[1066],seed[858],seed[1664],seed[290],seed[1475],seed[173],seed[593],seed[1700],seed[2329],seed[1479],seed[2902],seed[2476],seed[3190],seed[1370],seed[720],seed[70],seed[3810],seed[3984],seed[1313],seed[3903],seed[3684],seed[1832],seed[2138],seed[992],seed[1732],seed[2331],seed[2424],seed[3522],seed[3461],seed[1392],seed[1825],seed[14],seed[3837],seed[1647],seed[2719],seed[3973],seed[878],seed[1109],seed[3133],seed[2009],seed[1638],seed[1606],seed[3750],seed[3091],seed[4011],seed[22],seed[2217],seed[1938],seed[1156],seed[321],seed[3883],seed[274],seed[1788],seed[839],seed[500],seed[1054],seed[622],seed[3449],seed[558],seed[1979],seed[3196],seed[2198],seed[802],seed[2898],seed[2555],seed[3468],seed[2163],seed[2287],seed[2054],seed[3822],seed[380],seed[1798],seed[2783],seed[3019],seed[72],seed[2445],seed[1105],seed[913],seed[717],seed[79],seed[1472],seed[513],seed[753],seed[4073],seed[1355],seed[1764],seed[1219],seed[3334],seed[777],seed[1703],seed[3475],seed[1714],seed[2569],seed[2934],seed[3418],seed[1356],seed[2289],seed[1993],seed[1262],seed[218],seed[3452],seed[2239],seed[238],seed[2000],seed[134],seed[2829],seed[194],seed[3474],seed[1412],seed[2119],seed[2519],seed[3244],seed[3953],seed[1685],seed[387],seed[2602],seed[3399],seed[1780],seed[3902],seed[620],seed[4085],seed[1861],seed[2246],seed[3624],seed[7],seed[752],seed[3679],seed[3900],seed[3459],seed[1787],seed[1481],seed[2791],seed[1888],seed[772],seed[3456],seed[2200],seed[933],seed[3230],seed[3301],seed[3250],seed[638],seed[3650],seed[3165],seed[1252],seed[1341],seed[3185],seed[2270],seed[577],seed[75],seed[3228],seed[3321],seed[1395],seed[3266],seed[1801],seed[3048],seed[1199],seed[3239],seed[1722],seed[3577],seed[1797],seed[2658],seed[671],seed[3286],seed[2300],seed[543],seed[2276],seed[3129],seed[1433],seed[2525],seed[2982],seed[2883],seed[2177],seed[3588],seed[1741],seed[0],seed[2641],seed[711],seed[636],seed[3772],seed[1925],seed[11],seed[4084],seed[421],seed[2486],seed[1599],seed[3861],seed[3031],seed[1038],seed[936],seed[970],seed[1602],seed[1581],seed[1642],seed[1923],seed[1017],seed[2491],seed[3812],seed[954],seed[3834],seed[3023],seed[2110],seed[1070],seed[614],seed[226],seed[1235],seed[1237],seed[998],seed[3875],seed[2709],seed[272],seed[1662],seed[1418],seed[694],seed[2933],seed[3383],seed[1065],seed[3654],seed[2638],seed[1002],seed[1404],seed[3106],seed[2878],seed[2481],seed[2266],seed[3939],seed[3311],seed[91],seed[1646],seed[123],seed[3319],seed[346],seed[625],seed[1220],seed[3056],seed[552],seed[2520],seed[1608],seed[2976],seed[3741],seed[165],seed[2640],seed[2528],seed[2634],seed[849],seed[2670],seed[3170],seed[1360],seed[2745],seed[3534],seed[609],seed[2969],seed[1290],seed[334],seed[2739],seed[168],seed[1119],seed[1261],seed[4031],seed[2249],seed[3612],seed[2688],seed[3818],seed[2428],seed[1942],seed[1100],seed[32],seed[2694],seed[1128],seed[480],seed[1693],seed[1727],seed[1684],seed[606],seed[670],seed[1820],seed[2511],seed[1171],seed[3030],seed[3874],seed[974],seed[1879],seed[586],seed[214],seed[3663],seed[1434],seed[2241],seed[1476],seed[1603],seed[353],seed[197],seed[1030],seed[3672],seed[2070],seed[343],seed[3690],seed[776],seed[1342],seed[2553],seed[3860],seed[2433],seed[3993],seed[587],seed[3478],seed[3357],seed[3651],seed[983],seed[3674],seed[940],seed[3118],seed[2291],seed[1678],seed[1343],seed[3623],seed[3581],seed[385],seed[901],seed[1557],seed[1853],seed[3536],seed[3541],seed[835],seed[963],seed[966],seed[1967],seed[812],seed[3269],seed[3634],seed[3580],seed[2371],seed[3184],seed[1598],seed[3167],seed[1511],seed[2539],seed[328],seed[3192],seed[3070],seed[3508],seed[1755],seed[2611],seed[4018],seed[2388],seed[773],seed[3377],seed[3227],seed[3348],seed[3201],seed[2687],seed[3427],seed[1113],seed[3130],seed[642],seed[2037],seed[2697],seed[3896],seed[2404],seed[895],seed[1568],seed[828],seed[317],seed[607],seed[1738],seed[397],seed[185],seed[2112],seed[3374],seed[1743],seed[330],seed[3008],seed[121],seed[3120],seed[791],seed[1492],seed[146],seed[1391],seed[1966],seed[4070],seed[1203],seed[1924],seed[2209],seed[2190],seed[152],seed[1240],seed[427],seed[497],seed[2173],seed[2418],seed[4075],seed[1445],seed[1234],seed[1834],seed[3988],seed[2087],seed[490],seed[1450],seed[4074],seed[1566],seed[3142],seed[1502],seed[1828],seed[148],seed[3839],seed[600],seed[3929],seed[962],seed[659],seed[1477],seed[1175],seed[2204],seed[270],seed[2237],seed[323],seed[3096],seed[2164],seed[646],seed[3671],seed[257],seed[1707],seed[975],seed[626],seed[1332],seed[3174],seed[2873],seed[2800],seed[426],seed[2338],seed[1800],seed[2421],seed[2236],seed[2063],seed[1058],seed[3698],seed[3209],seed[544],seed[461],seed[2834],seed[1202],seed[2452],seed[3597],seed[2328],seed[3713],seed[1265],seed[3448],seed[326],seed[2129],seed[475],seed[3075],seed[655],seed[2517],seed[1486],seed[3670],seed[3846],seed[1555],seed[4043],seed[437],seed[483],seed[3972],seed[1032],seed[2534],seed[2787],seed[3497],seed[1056],seed[3708],seed[4009],seed[3119],seed[3290],seed[845],seed[2225],seed[925],seed[3969],seed[252],seed[3640],seed[2767],seed[3578],seed[3143],seed[3649],seed[889],seed[755],seed[3262],seed[2345],seed[589],seed[3287],seed[1806],seed[1372],seed[3783],seed[3510],seed[209],seed[186],seed[1982],seed[1921],seed[3800],seed[3952],seed[2166],seed[273],seed[3136],seed[3216],seed[3450],seed[1763],seed[2508],seed[2247],seed[2264],seed[1672],seed[1487],seed[792],seed[3806],seed[352],seed[1594],seed[2696],seed[3699],seed[703],seed[3694],seed[2228],seed[3760],seed[436],seed[1060],seed[3214],seed[1556],seed[2636],seed[892],seed[2590],seed[3298],seed[1345],seed[4034],seed[3393],seed[171],seed[258],seed[2605],seed[616],seed[95],seed[391],seed[3498],seed[3080],seed[1115],seed[4066],seed[381],seed[3916],seed[1120],seed[2626],seed[3409],seed[1044],seed[3529],seed[2771],seed[1158],seed[1193],seed[2633],seed[2103],seed[2630],seed[3221],seed[3155],seed[1726],seed[3005],seed[3],seed[1102],seed[3242],seed[2178],seed[3703],seed[1325],seed[3976],seed[3154],seed[1340],seed[2625],seed[2339],seed[999],seed[189],seed[651],seed[71],seed[245],seed[90],seed[3044],seed[2133],seed[3176],seed[1292],seed[1067],seed[3616],seed[3355],seed[204],seed[3163],seed[1903],seed[1242],seed[1552],seed[363],seed[997],seed[2033],seed[2732],seed[1166],seed[2443],seed[3573],seed[1563],seed[3887],seed[1104],seed[2826],seed[1571],seed[2531],seed[3705],seed[94],seed[1393],seed[803],seed[514],seed[2320],seed[1737],seed[2436],seed[192],seed[3455],seed[2454],seed[355],seed[3851],seed[3058],seed[1592],seed[668],seed[647],seed[2055],seed[1491],seed[18],seed[2124],seed[1936],seed[3364],seed[1735],seed[3539],seed[300],seed[1144],seed[3922],seed[35],seed[1695],seed[362],seed[2501],seed[2256],seed[1937],seed[268],seed[676],seed[1748],seed[3530],seed[1474],seed[3105],seed[3639],seed[2446],seed[1123],seed[3467],seed[1155],seed[3256],seed[181],seed[2784],seed[738],seed[2248],seed[1671],seed[61],seed[813],seed[1734],seed[725],seed[683],seed[3645],seed[2056],seed[3487],seed[2095],seed[2317],seed[769],seed[1901],seed[1885],seed[3501],seed[2915],seed[1835],seed[4012],seed[1742],seed[2001],seed[3280],seed[2414],seed[1597],seed[2507],seed[1217],seed[906],seed[1406],seed[3182],seed[950],seed[1992],seed[3625],seed[3779],seed[3442],seed[3098],seed[3787],seed[1333],seed[782],seed[2387],seed[3935],seed[681],seed[2691],seed[3283],seed[3384],seed[2559],seed[1306],seed[1271],seed[2262],seed[443],seed[2187],seed[978],seed[2774],seed[2156],seed[3210],seed[3292],seed[2724],seed[3372],seed[654],seed[3349],seed[3681],seed[1337],seed[1653],seed[1413],seed[1253],seed[3309],seed[3103],seed[1462],seed[360],seed[116],seed[4],seed[3350],seed[2897],seed[2945],seed[2524],seed[1444],seed[526],seed[377],seed[503],seed[2882],seed[1244],seed[2677],seed[3367],seed[3435],seed[2435],seed[458],seed[667],seed[2325],seed[1124],seed[1210],seed[1526],seed[2972],seed[2468],seed[447],seed[2399],seed[2530],seed[3949],seed[2254],seed[1362],seed[2913],seed[3833],seed[2509],seed[2682],seed[327],seed[1229],seed[1540],seed[1539],seed[2458],seed[2208],seed[145],seed[2144],seed[356],seed[2604],seed[3491],seed[1218],seed[2025],seed[1534],seed[3353],seed[2425],seed[179],seed[383],seed[432],seed[2226],seed[3460],seed[2066],seed[3248],seed[3064],seed[1024],seed[3961],seed[3425],seed[3730],seed[1681],seed[2741],seed[2942],seed[692],seed[3500],seed[2465],seed[3344],seed[1953],seed[1083],seed[3463],seed[3893],seed[1644],seed[2948],seed[2810],seed[3669],seed[2985],seed[3203],seed[3029],seed[1405],seed[2858],seed[3486],seed[1200],seed[1468],seed[3514],seed[931],seed[2849],seed[766],seed[3965],seed[535],seed[3441],seed[412],seed[2848],seed[3584],seed[3177],seed[474],seed[3808],seed[33],seed[3134],seed[876],seed[133],seed[3371],seed[3794],seed[1280],seed[3282],seed[3489],seed[3270],seed[2304],seed[2456],seed[1758],seed[3656],seed[2868],seed[1087]}),
        .cross_prob(cross_prob),
        .codeword(codeword2),
        .received(received2)
        );
        
    bsc bsc3(
        .clk(clk),
        .reset(reset),
        .seed({seed[1918],seed[524],seed[3736],seed[2813],seed[199],seed[1877],seed[299],seed[1459],seed[3365],seed[1019],seed[550],seed[1652],seed[1815],seed[3082],seed[2685],seed[1261],seed[2778],seed[269],seed[1253],seed[710],seed[1408],seed[506],seed[3304],seed[3540],seed[4075],seed[3862],seed[3824],seed[2929],seed[3322],seed[1474],seed[1719],seed[1929],seed[940],seed[1973],seed[3816],seed[2149],seed[725],seed[3755],seed[2172],seed[572],seed[408],seed[1939],seed[607],seed[1956],seed[2419],seed[1892],seed[2129],seed[2101],seed[1917],seed[3835],seed[3552],seed[1433],seed[1429],seed[1205],seed[1716],seed[2193],seed[2287],seed[3668],seed[4050],seed[3993],seed[2092],seed[1188],seed[544],seed[585],seed[2808],seed[3687],seed[1507],seed[641],seed[1916],seed[2469],seed[2726],seed[3726],seed[1197],seed[3228],seed[870],seed[3520],seed[1931],seed[3600],seed[2661],seed[2875],seed[2632],seed[2576],seed[3371],seed[1386],seed[3264],seed[63],seed[1338],seed[2128],seed[1496],seed[1828],seed[2691],seed[2373],seed[221],seed[952],seed[4048],seed[4044],seed[289],seed[3339],seed[1935],seed[1388],seed[2806],seed[189],seed[875],seed[4014],seed[447],seed[336],seed[1802],seed[2209],seed[384],seed[1218],seed[2985],seed[3451],seed[1641],seed[169],seed[1219],seed[1048],seed[1660],seed[713],seed[2820],seed[201],seed[3970],seed[1453],seed[1961],seed[1899],seed[1689],seed[3751],seed[2647],seed[900],seed[2842],seed[3455],seed[3899],seed[3914],seed[3605],seed[1572],seed[1708],seed[1469],seed[172],seed[3599],seed[37],seed[2038],seed[1791],seed[1749],seed[87],seed[1411],seed[2925],seed[1810],seed[2178],seed[534],seed[559],seed[1413],seed[2219],seed[1770],seed[797],seed[1982],seed[1706],seed[1595],seed[1705],seed[3399],seed[3139],seed[520],seed[3284],seed[1694],seed[3386],seed[565],seed[2447],seed[1299],seed[2829],seed[3793],seed[3700],seed[2918],seed[946],seed[3472],seed[1430],seed[2708],seed[3784],seed[263],seed[1883],seed[3693],seed[2672],seed[3996],seed[1552],seed[2170],seed[2237],seed[3646],seed[1966],seed[3643],seed[795],seed[1486],seed[1500],seed[467],seed[344],seed[1070],seed[3978],seed[3189],seed[3468],seed[2010],seed[3044],seed[2114],seed[3525],seed[1331],seed[3799],seed[1896],seed[3030],seed[4000],seed[3895],seed[3249],seed[883],seed[2700],seed[3613],seed[101],seed[1067],seed[3321],seed[874],seed[910],seed[2338],seed[2014],seed[3579],seed[1290],seed[3880],seed[906],seed[4043],seed[3967],seed[1281],seed[3834],seed[3923],seed[3063],seed[951],seed[2159],seed[1396],seed[1133],seed[329],seed[2322],seed[2750],seed[3195],seed[3889],seed[461],seed[3596],seed[2906],seed[3194],seed[1954],seed[3663],seed[3572],seed[1034],seed[1189],seed[2874],seed[3220],seed[53],seed[3795],seed[3533],seed[2481],seed[1844],seed[3404],seed[1318],seed[876],seed[3725],seed[639],seed[3919],seed[1087],seed[1555],seed[3803],seed[3577],seed[688],seed[2033],seed[3670],seed[2723],seed[2527],seed[786],seed[3746],seed[3181],seed[2085],seed[827],seed[2274],seed[1225],seed[4045],seed[252],seed[848],seed[1995],seed[2939],seed[94],seed[2834],seed[2735],seed[3580],seed[707],seed[1293],seed[3872],seed[2069],seed[2586],seed[1107],seed[3252],seed[1126],seed[3944],seed[2956],seed[208],seed[4025],seed[3973],seed[2095],seed[1049],seed[370],seed[3820],seed[3684],seed[1646],seed[2553],seed[2658],seed[122],seed[2137],seed[110],seed[148],seed[250],seed[3230],seed[2998],seed[1680],seed[1728],seed[3639],seed[1406],seed[1339],seed[3283],seed[3175],seed[1403],seed[4076],seed[1276],seed[2291],seed[2724],seed[987],seed[790],seed[1981],seed[484],seed[308],seed[1970],seed[2690],seed[115],seed[2627],seed[3591],seed[950],seed[2961],seed[989],seed[1251],seed[3859],seed[1380],seed[3361],seed[3214],seed[2802],seed[3825],seed[3818],seed[2540],seed[1834],seed[3086],seed[3901],seed[594],seed[1351],seed[3109],seed[2649],seed[1059],seed[1332],seed[2432],seed[4091],seed[2221],seed[1540],seed[497],seed[43],seed[3417],seed[1950],seed[2043],seed[3062],seed[420],seed[1495],seed[567],seed[712],seed[2631],seed[1946],seed[1988],seed[2940],seed[1588],seed[3033],seed[1300],seed[752],seed[3936],seed[1013],seed[316],seed[1710],seed[1359],seed[369],seed[3647],seed[2602],seed[1852],seed[1887],seed[2339],seed[2155],seed[3683],seed[3458],seed[1608],seed[3958],seed[4090],seed[719],seed[241],seed[501],seed[1817],seed[3087],seed[185],seed[2119],seed[3509],seed[2],seed[652],seed[3383],seed[2941],seed[2667],seed[2390],seed[2046],seed[1944],seed[2548],seed[3966],seed[3989],seed[2427],seed[334],seed[637],seed[1444],seed[3065],seed[2888],seed[3446],seed[967],seed[2426],seed[3499],seed[3794],seed[2465],seed[3199],seed[574],seed[805],seed[2721],seed[311],seed[895],seed[464],seed[2276],seed[3396],seed[616],seed[3720],seed[3701],seed[538],seed[3301],seed[3166],seed[3257],seed[3131],seed[1236],seed[3573],seed[1229],seed[1230],seed[291],seed[2972],seed[2747],seed[292],seed[1745],seed[3001],seed[2135],seed[4006],seed[1357],seed[1704],seed[3436],seed[1523],seed[728],seed[1957],seed[1363],seed[1120],seed[1860],seed[4060],seed[1836],seed[1135],seed[1978],seed[1057],seed[621],seed[2551],seed[2230],seed[2899],seed[166],seed[1132],seed[936],seed[2120],seed[4047],seed[3717],seed[2962],seed[1266],seed[4092],seed[434],seed[1687],seed[3928],seed[2526],seed[3084],seed[379],seed[1161],seed[153],seed[4023],seed[774],seed[1930],seed[1894],seed[3187],seed[824],seed[1167],seed[3739],seed[1345],seed[2652],seed[3129],seed[1808],seed[74],seed[1594],seed[2454],seed[1385],seed[2885],seed[3539],seed[2964],seed[3753],seed[3363],seed[999],seed[1115],seed[38],seed[3459],seed[566],seed[2588],seed[2388],seed[1675],seed[3992],seed[1833],seed[1228],seed[1162],seed[2883],seed[1454],seed[2959],seed[1378],seed[3542],seed[3984],seed[1438],seed[2694],seed[318],seed[2025],seed[2444],seed[1280],seed[401],seed[3735],seed[613],seed[3756],seed[3217],seed[2760],seed[1233],seed[1481],seed[664],seed[2289],seed[3903],seed[2688],seed[3118],seed[3096],seed[3508],seed[1574],seed[2541],seed[1211],seed[1042],seed[2977],seed[3790],seed[3535],seed[481],seed[4008],seed[3526],seed[894],seed[3348],seed[1150],seed[3607],seed[1907],seed[1798],seed[2657],seed[3057],seed[88],seed[2697],seed[2379],seed[846],seed[1461],seed[954],seed[1544],seed[1451],seed[322],seed[355],seed[3406],seed[61],seed[210],seed[3122],seed[246],seed[2232],seed[2845],seed[2366],seed[2107],seed[3275],seed[541],seed[1110],seed[3527],seed[1457],seed[599],seed[3940],seed[3211],seed[701],seed[1392],seed[3886],seed[2909],seed[368],seed[3904],seed[2130],seed[182],seed[643],seed[2668],seed[3776],seed[2116],seed[1854],seed[96],seed[1789],seed[2403],seed[662],seed[1005],seed[2325],seed[400],seed[422],seed[2318],seed[1144],seed[1835],seed[2425],seed[3051],seed[2570],seed[2686],seed[3185],seed[3948],seed[3715],seed[3203],seed[2531],seed[1482],seed[1171],seed[86],seed[1399],seed[347],seed[124],seed[2800],seed[1725],seed[610],seed[3495],seed[290],seed[2635],seed[360],seed[2392],seed[78],seed[3375],seed[403],seed[2236],seed[3298],seed[4069],seed[2568],seed[2642],seed[1605],seed[3208],seed[668],seed[959],seed[2436],seed[3402],seed[186],seed[2995],seed[2293],seed[2294],seed[684],seed[1627],seed[3467],seed[2645],seed[3937],seed[2249],seed[321],seed[1764],seed[3150],seed[2393],seed[986],seed[1170],seed[2204],seed[1124],seed[3713],seed[3961],seed[1222],seed[3877],seed[2771],seed[676],seed[3870],seed[1422],seed[1562],seed[2165],seed[1784],seed[1800],seed[2943],seed[1296],seed[2422],seed[1409],seed[1452],seed[980],seed[1591],seed[1759],seed[861],seed[976],seed[2220],seed[33],seed[551],seed[1510],seed[1941],seed[2613],seed[3170],seed[146],seed[3100],seed[2559],seed[3123],seed[2766],seed[1282],seed[2917],seed[3390],seed[1576],seed[1185],seed[3113],seed[3716],seed[242],seed[2870],seed[3570],seed[2539],seed[4061],seed[3832],seed[837],seed[3661],seed[3916],seed[77],seed[1558],seed[305],seed[3077],seed[1116],seed[3318],seed[2983],seed[1794],seed[2757],seed[530],seed[3069],seed[836],seed[82],seed[2718],seed[1658],seed[2256],seed[111],seed[294],seed[1095],seed[2493],seed[781],seed[2184],seed[1928],seed[3838],seed[3445],seed[132],seed[812],seed[228],seed[1766],seed[921],seed[2597],seed[1182],seed[759],seed[2081],seed[964],seed[2630],seed[3733],seed[2612],seed[720],seed[1414],seed[2516],seed[3],seed[1682],seed[2368],seed[2039],seed[3632],seed[508],seed[2653],seed[2810],seed[1543],seed[2618],seed[3091],seed[2121],seed[922],seed[1448],seed[19],seed[2138],seed[1865],seed[239],seed[1200],seed[1043],seed[2755],seed[313],seed[2185],seed[1033],seed[691],seed[1686],seed[2409],seed[1653],seed[2126],seed[3206],seed[1440],seed[1202],seed[1746],seed[771],seed[4004],seed[2850],seed[222],seed[855],seed[3863],seed[3188],seed[2664],seed[1934],seed[3556],seed[1948],seed[636],seed[1097],seed[3202],seed[2903],seed[3602],seed[2103],seed[3688],seed[2681],seed[2737],seed[2509],seed[2495],seed[681],seed[6],seed[4066],seed[1822],seed[3681],seed[1436],seed[3637],seed[1437],seed[2946],seed[387],seed[730],seed[2206],seed[801],seed[474],seed[2327],seed[1164],seed[653],seed[2824],seed[2313],seed[3629],seed[978],seed[1714],seed[273],seed[749],seed[1733],seed[1175],seed[1547],seed[341],seed[2163],seed[348],seed[3172],seed[1991],seed[1602],seed[1137],seed[2110],seed[949],seed[808],seed[90],seed[3289],seed[2633],seed[3812],seed[340],seed[2926],seed[2024],seed[1927],seed[528],seed[3169],seed[4080],seed[804],seed[984],seed[729],seed[1141],seed[3448],seed[2317],seed[3505],seed[1569],seed[13],seed[1294],seed[825],seed[1659],seed[1855],seed[3900],seed[3317],seed[3089],seed[2817],seed[3822],seed[2836],seed[1045],seed[69],seed[3503],seed[3939],seed[3486],seed[1925],seed[2467],seed[1681],seed[1509],seed[1308],seed[2355],seed[452],seed[2462],seed[939],seed[1484],seed[3890],seed[1631],seed[3878],seed[767],seed[1751],seed[2345],seed[2933],seed[857],seed[934],seed[1153],seed[2947],seed[919],seed[410],seed[3130],seed[1151],seed[1667],seed[2975],seed[3652],seed[397],seed[31],seed[2458],seed[207],seed[3792],seed[3360],seed[3142],seed[3098],seed[3487],seed[2648],seed[3039],seed[1581],seed[438],seed[1499],seed[3453],seed[2329],seed[1888],seed[2854],seed[1169],seed[658],seed[1012],seed[439],seed[1367],seed[615],seed[2756],seed[2186],seed[1405],seed[376],seed[1063],seed[3427],seed[3623],seed[2793],seed[2019],seed[3857],seed[256],seed[671],seed[3247],seed[489],seed[892],seed[2240],seed[2616],seed[3915],seed[2871],seed[249],seed[3584],seed[3023],seed[3490],seed[1748],seed[721],seed[1753],seed[1598],seed[2394],seed[247],seed[2582],seed[3676],seed[365],seed[3034],seed[2740],seed[2535],seed[2518],seed[2448],seed[1382],seed[2063],seed[3235],seed[1297],seed[300],seed[204],seed[2260],seed[298],seed[3461],seed[114],seed[3642],seed[3828],seed[2936],seed[3551],seed[2594],seed[920],seed[1341],seed[1636],seed[2188],seed[4084],seed[1769],seed[1479],seed[3771],seed[1721],seed[4019],seed[1435],seed[1609],seed[2573],seed[2980],seed[1584],seed[1573],seed[3737],seed[4028],seed[1096],seed[3002],seed[457],seed[3036],seed[1007],seed[3485],seed[3645],seed[42],seed[2158],seed[3013],seed[3773],seed[1289],seed[811],seed[692],seed[58],seed[1214],seed[3968],seed[2336],seed[3450],seed[2018],seed[2272],seed[2124],seed[1355],seed[8],seed[822],seed[445],seed[3982],seed[319],seed[3059],seed[359],seed[1303],seed[1804],seed[2670],seed[2361],seed[3950],seed[64],seed[3601],seed[320],seed[1314],seed[1123],seed[869],seed[1023],seed[3161],seed[2791],seed[2468],seed[1513],seed[2797],seed[3778],seed[1824],seed[1203],seed[2253],seed[2769],seed[3581],seed[1768],seed[212],seed[3070],seed[1799],seed[3243],seed[193],seed[1397],seed[3180],seed[2752],seed[3549],seed[1945],seed[1638],seed[871],seed[2510],seed[682],seed[2026],seed[3764],seed[2442],seed[3927],seed[898],seed[2433],seed[120],seed[2315],seed[1893],seed[3798],seed[2604],seed[3564],seed[4052],seed[1348],seed[3852],seed[2037],seed[3336],seed[1320],seed[1747],seed[1587],seed[849],seed[1718],seed[2877],seed[1691],seed[3014],seed[3842],seed[1585],seed[3456],seed[192],seed[555],seed[753],seed[765],seed[744],seed[460],seed[2146],seed[1617],seed[638],seed[624],seed[2900],seed[2279],seed[3567],seed[34],seed[3072],seed[1736],seed[1535],seed[2528],seed[3775],seed[3053],seed[1254],seed[2584],seed[1343],seed[1017],seed[2581],seed[3562],seed[1387],seed[2087],seed[2572],seed[349],seed[473],seed[1467],seed[1616],seed[665],seed[2734],seed[4071],seed[3484],seed[151],seed[1996],seed[3644],seed[1078],seed[659],seed[2957],seed[3806],seed[2380],seed[202],seed[2713],seed[3494],seed[2567],seed[93],seed[686],seed[2628],seed[3514],seed[3251],seed[1058],seed[1897],seed[179],seed[2153],seed[2781],seed[2286],seed[3530],seed[740],seed[1779],seed[2994],seed[3752],seed[4081],seed[2898],seed[3449],seed[1027],seed[2076],seed[620],seed[3327],seed[1093],seed[138],seed[3424],seed[3209],seed[2514],seed[2763],seed[1047],seed[2464],seed[2320],seed[3610],seed[1538],seed[913],seed[1490],seed[2910],seed[3938],seed[3625],seed[450],seed[66],seed[3388],seed[236],seed[2984],seed[618],seed[1503],seed[449],seed[2342],seed[332],seed[220],seed[799],seed[3976],seed[2938],seed[4085],seed[4005],seed[750],seed[3179],seed[29],seed[2408],seed[3239],seed[2908],seed[1674],seed[310],seed[2386],seed[2140],seed[3529],seed[902],seed[864],seed[2682],seed[3922],seed[2494],seed[3302],seed[2415],seed[1878],seed[3557],seed[1416],seed[3658],seed[2471],seed[1163],seed[2118],seed[703],seed[1801],seed[1599],seed[3628],seed[1709],seed[1642],seed[928],seed[539],seed[1909],seed[3429],seed[1589],seed[3991],seed[2125],seed[806],seed[1391],seed[312],seed[2387],seed[1879],seed[2477],seed[134],seed[1084],seed[1707],seed[2349],seed[3924],seed[363],seed[3350],seed[3391],seed[2154],seed[492],seed[331],seed[2203],seed[1053],seed[1847],seed[1781],seed[1821],seed[2405],seed[361],seed[2347],seed[971],seed[3151],seed[2323],seed[2078],seed[260],seed[3121],seed[4030],seed[3972],seed[2701],seed[1895],seed[1076],seed[1298],seed[4059],seed[882],seed[118],seed[1842],seed[2189],seed[3691],seed[1625],seed[76],seed[3589],seed[4073],seed[1761],seed[398],seed[1172],seed[3860],seed[562],seed[431],seed[852],seed[2575],seed[746],seed[3699],seed[1943],seed[1669],seed[3017],seed[4031],seed[3430],seed[1088],seed[1178],seed[2190],seed[1863],seed[796],seed[1313],seed[1536],seed[858],seed[2466],seed[3821],seed[328],seed[2952],seed[516],seed[1183],seed[1323],seed[2622],seed[3074],seed[1922],seed[2549],seed[2222],seed[2143],seed[1592],seed[549],seed[3782],seed[2480],seed[2695],seed[3810],seed[2171],seed[3167],seed[2304],seed[3867],seed[3473],seed[788],seed[927],seed[3758],seed[2546],seed[2953],seed[3101],seed[1551],seed[3364],seed[2765],seed[1149],seed[838],seed[741],seed[28],seed[2876],seed[3474],seed[3411],seed[2057],seed[2067],seed[649],seed[734],seed[859],seed[3910],seed[2428],seed[3042],seed[1156],seed[2297],seed[3695],seed[2678],seed[1243],seed[200],seed[3397],seed[3774],seed[3696],seed[2707],seed[695],seed[1340],seed[1977],seed[2683],seed[377],seed[3447],seed[24],seed[1903],seed[3270],seed[3897],seed[209],seed[3442],seed[509],seed[2201],seed[3431],seed[2319],seed[885],seed[3544],seed[302],seed[630],seed[2932],seed[3041],seed[582],seed[3518],seed[218],seed[1241],seed[3127],seed[2866],seed[2267],seed[1419],seed[1038],seed[3560],seed[556],seed[2865],seed[2732],seed[68],seed[1514],seed[1008],seed[1328],seed[1870],seed[1002],seed[4032],seed[1985],seed[1864],seed[1624],seed[650],seed[338],seed[2555],seed[798],seed[2981],seed[2239],seed[909],seed[1545],seed[3236],seed[1434],seed[2020],seed[1035],seed[1557],seed[140],seed[3193],seed[2215],seed[961],seed[1142],seed[2282],seed[3787],seed[1426],seed[2591],seed[1011],seed[1740],seed[2410],seed[3231],seed[2411],seed[500],seed[2071],seed[3802],seed[2423],seed[1213],seed[433],seed[4013],seed[1094],seed[2292],seed[1356],seed[1867],seed[972],seed[3744],seed[850],seed[561],seed[3040],seed[3480],seed[742],seed[1190],seed[1868],seed[3233],seed[1906],seed[2086],seed[3745],seed[2229],seed[589],seed[933],seed[2132],seed[1064],seed[1085],seed[3067],seed[2809],seed[2441],seed[1654],seed[2950],seed[123],seed[1069],seed[3392],seed[1517],seed[1117],seed[3921],seed[1738],seed[1611],seed[133],seed[2619],seed[416],seed[3957],seed[1990],seed[3528],seed[1676],seed[2934],seed[2725],seed[3465],seed[1317],seed[493],seed[1677],seed[2461],seed[1284],seed[2285],seed[3641],seed[3705],seed[3075],seed[2788],seed[307],seed[3104],seed[2102],seed[14],seed[3163],seed[35],seed[2601],seed[3140],seed[3594],seed[174],seed[2484],seed[2916],seed[2307],seed[1607],seed[4036],seed[1130],seed[685],seed[3258],seed[3242],seed[119],seed[1793],seed[2060],seed[3561],seed[2712],seed[285],seed[2202],seed[2692],seed[2169],seed[3734],seed[2115],seed[3523],seed[2271],seed[4058],seed[1932],seed[581],seed[2758],seed[3708],seed[2585],seed[1335],seed[3826],seed[2547],seed[1744],seed[3489],seed[1637],seed[2344],seed[257],seed[3638],seed[2736],seed[3421],seed[1809],seed[1104],seed[2492],seed[2055],seed[3656],seed[1373],seed[588],seed[155],seed[1431],seed[1001],seed[2098],seed[3657],seed[107],seed[458],seed[2151],seed[1065],seed[57],seed[230],seed[205],seed[337],seed[40],seed[823],seed[1610],seed[1987],seed[2174],seed[1622],seed[167],seed[2210],seed[1623],seed[514],seed[1797],seed[595],seed[3016],seed[1267],seed[675],seed[648],seed[1737],seed[2655],seed[1106],seed[3918],seed[2892],seed[994],seed[1603],seed[3439],seed[2574],seed[3614],seed[3955],seed[2663],seed[975],seed[326],seed[758],seed[2283],seed[644],seed[2669],seed[766],seed[3454],seed[1796],seed[2389],seed[3300],seed[109],seed[3830],seed[814],seed[737],seed[2414],seed[2181],seed[3291],seed[1811],seed[2895],seed[718],seed[1711],seed[2812],seed[2679],seed[2557],seed[2993],seed[3340],seed[1285],seed[4093],seed[2047],seed[1235],seed[52],seed[2162],seed[3315],seed[2248],seed[2131],seed[258],seed[3931],seed[723],seed[3401],seed[3722],seed[26],seed[3709],seed[3149],seed[2006],seed[2935],seed[3056],seed[918],seed[2930],seed[633],seed[3460],seed[1920],seed[465],seed[2911],seed[2945],seed[2073],seed[5],seed[2455],seed[12],seed[1566],seed[698],seed[3960],seed[1309],seed[1006],seed[3341],seed[2357],seed[754],seed[3788],seed[2571],seed[1635],seed[2569],seed[195],seed[2815],seed[1720],seed[3706],seed[619],seed[288],seed[2218],seed[1492],seed[1952],seed[942],seed[3428],seed[1274],seed[1805],seed[270],seed[27],seed[3945],seed[444],seed[2328],seed[1021],seed[3515],seed[896],seed[309],seed[1644],seed[1795],seed[3779],seed[3232],seed[3409],seed[54],seed[1127],seed[494],seed[10],seed[571],seed[1840],seed[2879],seed[1614],seed[3005],seed[383],seed[2000],seed[352],seed[745],seed[944],seed[3225],seed[2988],seed[1307],seed[2774],seed[411],seed[1861],seed[1501],seed[904],seed[2564],seed[345],seed[2008],seed[2790],seed[1292],seed[1354],seed[2714],seed[1061],seed[583],seed[2792],seed[2265],seed[3332],seed[1962],seed[2262],seed[3178],seed[1372],seed[3124],seed[1083],seed[3303],seed[1288],seed[3833],seed[1152],seed[860],seed[275],seed[4018],seed[2651],seed[2644],seed[1633],seed[731],seed[213],seed[960],seed[2301],seed[3664],seed[1882],seed[793],seed[2872],seed[2122],seed[2108],seed[791],seed[2522],seed[3959],seed[3215],seed[2491],seed[3478],seed[3061],seed[2275],seed[59],seed[1287],seed[3675],seed[1109],seed[3543],seed[1324],seed[2023],seed[1712],seed[2029],seed[1091],seed[1407],seed[1498],seed[780],seed[2521],seed[1112],seed[2704],seed[3221],seed[1086],seed[1819],seed[3168],seed[907],seed[440],seed[1643],seed[2828],seed[611],seed[2051],seed[2263],seed[157],seed[3854],seed[1814],seed[3165],seed[1512],seed[1221],seed[3492],seed[1938],seed[2015],seed[789],seed[462],seed[3712],seed[3855],seed[1488],seed[1337],seed[569],seed[702],seed[2992],seed[0],seed[779],seed[3980],seed[164],seed[1301],seed[446],seed[1724],seed[3319],seed[2727],seed[511],seed[2839],seed[635],seed[1757],seed[603],seed[3634],seed[3942],seed[2430],seed[2331],seed[552],seed[3006],seed[1333],seed[2213],seed[2767],seed[518],seed[393],seed[3772],seed[667],seed[2924],seed[1729],seed[2278],seed[3356],seed[394],seed[1302],seed[3585],seed[196],seed[2578],seed[1255],seed[2280],seed[1304],seed[2333],seed[39],seed[3156],seed[2748],seed[997],seed[2214],seed[362],seed[844],seed[3240],seed[1311],seed[2673],seed[602],seed[2109],seed[1483],seed[1726],seed[1739],seed[3387],seed[343],seed[2965],seed[1291],seed[1604],seed[2951],seed[2354],seed[3612],seed[2141],seed[1959],seed[598],seed[3441],seed[2486],seed[1071],seed[3471],seed[2375],seed[2852],seed[1976],seed[1975],seed[1765],seed[1319],seed[3229],seed[1730],seed[1525],seed[2884],seed[3144],seed[3320],seed[3182],seed[3254],seed[628],seed[1381],seed[998],seed[2923],seed[1553],seed[1734],seed[899],seed[1515],seed[2978],seed[935],seed[760],seed[1942],seed[206],seed[925],seed[2247],seed[2782],seed[3433],seed[1018],seed[1619],seed[3029],seed[2134],seed[3164],seed[819],seed[2543],seed[265],seed[2580],seed[2050],seed[3135],seed[2905],seed[672],seed[1275],seed[18],seed[802],seed[716],seed[188],seed[223],seed[2352],seed[3674],seed[2383],seed[3907],seed[264],seed[3650],seed[2634],seed[1816],seed[3537],seed[3975],seed[3714],seed[4042],seed[1108],seed[2284],seed[1030],seed[105],seed[3218],seed[1493],seed[2300],seed[3609],seed[480],seed[1648],seed[346],seed[3197],seed[577],seed[2053],seed[3212],seed[924],seed[3060],seed[1655],seed[2893],seed[938],seed[79],seed[1081],seed[3358],seed[44],seed[2759],seed[131],seed[3586],seed[1477],seed[2840],seed[3868],seed[1803],seed[1400],seed[1999],seed[1541],seed[2048],seed[2646],seed[2034],seed[4002],seed[3250],seed[1259],seed[2517],seed[1516],seed[3416],seed[2452],seed[2127],seed[3483],seed[3626],seed[3479],seed[2823],seed[2266],seed[3248],seed[2459],seed[903],seed[1364],seed[1993],seed[3545],seed[3031],seed[2927],seed[325],seed[2536],seed[1231],seed[623],seed[415],seed[2017],seed[226],seed[3049],seed[2070],seed[219],seed[3425],seed[663],seed[2963],seed[2662],seed[564],seed[1402],seed[2420],seed[3045],seed[4034],seed[1365],seed[3174],seed[1664],seed[2506],seed[1080],seed[3521],seed[3353],seed[1131],seed[1914],seed[1068],seed[533],seed[1837],seed[1195],seed[3011],seed[884],seed[3400],seed[2890],seed[3690],seed[3136],seed[722],seed[3234],seed[3080],seed[1249],seed[2579],seed[977],seed[2715],seed[1665],seed[3437],seed[3702],seed[3742],seed[3731],seed[1898],seed[3692],seed[2948],seed[425],seed[3963],seed[979],seed[2161],seed[1165],seed[2052],seed[738],seed[1508],seed[3905],seed[600],seed[1915],seed[2478],seed[2443],seed[194],seed[1783],seed[3423],seed[1891],seed[1208],seed[259],seed[1196],seed[632],seed[1874],seed[380],seed[834],seed[2913],seed[3097],seed[2299],seed[3032],seed[2717],seed[11],seed[2421],seed[1632],seed[1775],seed[48],seed[2534],seed[1077],seed[1849],seed[3078],seed[1758],seed[3463],seed[1550],seed[553],seed[2861],seed[1082],seed[3438],seed[2321],seed[3226],seed[3892],seed[423],seed[2489],seed[2650],seed[2111],seed[2356],seed[2860],seed[2439],seed[974],seed[3493],seed[1024],seed[2722],seed[957],seed[3906],seed[3883],seed[1401],seed[3162],seed[1210],seed[2970],seed[1786],seed[941],seed[3920],seed[382],seed[3384],seed[2639],seed[1447],seed[3488],seed[626],seed[2314],seed[2805],seed[521],seed[2955],seed[1851],seed[3583],seed[1556],seed[726],seed[3640],seed[102],seed[1671],seed[2991],seed[2787],seed[931],seed[1232],seed[1806],seed[2529],seed[2498],seed[1839],seed[356],seed[2835],seed[1342],seed[476],seed[3286],seed[3055],seed[3929],seed[646],seed[95],seed[2113],seed[1845],seed[592],seed[1040],seed[841],seed[3134],seed[3048],seed[262],seed[908],seed[315],seed[2058],seed[1848],seed[593],seed[3237],seed[141],seed[1666],seed[3593],seed[3146],seed[3207],seed[631],seed[3079],seed[2391],seed[459],seed[1923],seed[3050],seed[3721],seed[3590],seed[1546],seed[3947],seed[1924],seed[498],seed[654],seed[277],seed[1717],seed[130],seed[2878],seed[968],seed[1468],seed[1240],seed[2838],seed[2590],seed[1125],seed[2777],seed[3845],seed[1394],seed[2511],seed[171],seed[2507],seed[914],seed[1020],seed[22],seed[388],seed[622],seed[49],seed[1846],seed[2479],seed[661],seed[724],seed[576],seed[266],seed[211],seed[579],seed[1361],seed[3395],seed[818],seed[2659],seed[2360],seed[2742],seed[1843],seed[1174],seed[296],seed[2770],seed[3724],seed[424],seed[2561],seed[1537],seed[1480],seed[981],seed[3550],seed[1969],seed[2921],seed[1412],seed[3502],seed[2841],seed[32],seed[2979],seed[2160],seed[1963],seed[3081],seed[3669],seed[2680],seed[3273],seed[1039],seed[1439],seed[1277],seed[2621],seed[873],seed[330],seed[1606],seed[2346],seed[3770],seed[2485],seed[3342],seed[2699],seed[4088],seed[2819],seed[178],seed[1528],seed[297],seed[3913],seed[647],seed[813],seed[4016],seed[1820],seed[2021],seed[3723],seed[3979],seed[3869],seed[170],seed[761],seed[863],seed[609],seed[2780],seed[3760],seed[1697],seed[342],seed[2863],seed[2001],seed[3804],seed[3111],seed[1158],seed[1960],seed[286],seed[1022],seed[3470],seed[700],seed[1441],seed[3413],seed[1857],seed[1889],seed[472],seed[1875],seed[2090],seed[2156],seed[679],seed[2487],seed[1521],seed[1148],seed[3815],seed[3732],seed[3635],seed[317],seed[830],seed[777],seed[504],seed[406],seed[1360],seed[739],seed[608],seed[3500],seed[1983],seed[2112],seed[2603],seed[2363],seed[512],seed[792],seed[432],seed[3837],seed[3279],seed[2552],seed[1118],seed[563],seed[3861],seed[3743],seed[85],seed[1613],seed[2512],seed[2144],seed[3685],seed[244],seed[546],seed[2438],seed[1398],seed[666],seed[1262],seed[3326],seed[2460],seed[165],seed[1621],seed[2105],seed[3337],seed[4024],seed[2503],seed[3578],seed[231],seed[1187],seed[3466],seed[2896],seed[3263],seed[3819],seed[1050],seed[333],seed[655],seed[3147],seed[3280],seed[2869],seed[1004],seed[3783],seed[4027],seed[3686],seed[3757],seed[2577],seed[2281],seed[3874],seed[2164],seed[2372],seed[3064],seed[97],seed[485],seed[2675],seed[851],seed[3844],seed[2225],seed[2592],seed[3654],seed[2401],seed[2505],seed[1559],seed[1286],seed[1979],seed[1143],seed[4077],seed[1154],seed[3606],seed[98],seed[3378],seed[3698],seed[2523],seed[1194],seed[763],seed[502],seed[1168],seed[2196],seed[1217],seed[1044],seed[2728],seed[3849],seed[3035],seed[1271],seed[1458],seed[2607],seed[36],seed[2407],seed[25],seed[2967],seed[2335],seed[2402],seed[1994],seed[3491],seed[1329],seed[1445],seed[3673],seed[3276],seed[4003],seed[1463],seed[1651],seed[350],seed[2406],seed[2440],seed[278],seed[1869],seed[2180],seed[3374],seed[727],seed[390],seed[1443],seed[1756],seed[3865],seed[3009],seed[468],seed[2605],seed[1016],seed[1427],seed[3964],seed[1327],seed[229],seed[3046],seed[2711],seed[3323],seed[1206],seed[1368],seed[3718],seed[3205],seed[1701],seed[1511],seed[2273],seed[245],seed[2986],seed[3346],seed[966],seed[2326],seed[2937],seed[1121],seed[2175],seed[2072],seed[2623],seed[3912],seed[1974],seed[683],seed[3157],seed[1936],seed[15],seed[2099],seed[2542],seed[1578],seed[191],seed[690],seed[2233],seed[2949],seed[3324],seed[956],seed[2257],seed[251],seed[2041],seed[1529],seed[1138],seed[4049],seed[2397],seed[2049],seed[893],seed[816],seed[238],seed[3971],seed[2987],seed[1315],seed[3148],seed[2556],seed[62],seed[1224],seed[2768],seed[2028],seed[2011],seed[1829],seed[1777],seed[280],seed[3385],seed[2942],seed[3648],seed[3309],seed[3563],seed[287],seed[396],seed[1727],seed[2643],seed[3373],seed[2508],seed[2194],seed[3587],seed[807],seed[443],seed[2261],seed[2089],seed[1395],seed[113],seed[3022],seed[1014],seed[3848],seed[2902],seed[3740],seed[527],seed[399],seed[3133],seed[2996],seed[2207],seed[1989],seed[3008],seed[697],seed[3839],seed[2598],seed[1580],seed[2786],seed[926],seed[2083],seed[3297],seed[2901],seed[3112],seed[142],seed[748],seed[2565],seed[568],seed[601],seed[2334],seed[2826],seed[3797],seed[4021],seed[3224],seed[1628],seed[2859],seed[2123],seed[3253],seed[3555],seed[2997],seed[1812],seed[1940],seed[421],seed[2744],seed[3840],seed[536],seed[2032],seed[3926],seed[3325],seed[2147],seed[2068],seed[696],seed[2851],seed[711],seed[3271],seed[451],seed[1871],seed[3769],seed[1257],seed[1933],seed[1362],seed[3565],seed[3592],seed[2104],seed[366],seed[3719],seed[373],seed[3780],seed[2496],seed[2638],seed[1223],seed[1683],seed[2482],seed[3186],seed[670],seed[454],seed[1560],seed[1201],seed[143],seed[2016],seed[542],seed[535],seed[2928],seed[1539],seed[958],seed[4039],seed[1593],seed[854],seed[1237],seed[1446],seed[845],seed[2044],seed[1244],seed[1853],seed[1478],seed[3536],seed[2764],seed[3697],seed[3177],seed[303],seed[3246],seed[2666],seed[2803],seed[3120],seed[3138],seed[463],seed[435],seed[3043],seed[674],seed[3891],seed[1561],seed[4035],seed[1442],seed[2502],seed[3094],seed[3210],seed[831],seed[3888],seed[2295],seed[558],seed[3941],seed[3126],seed[1542],seed[2629],seed[3310],seed[2195],seed[1565],seed[1432],seed[83],seed[116],seed[3443],seed[3379],seed[2369],seed[3152],seed[1114],seed[1866],seed[3352],seed[879],seed[2973],seed[800],seed[4087],seed[2676],seed[1713],seed[2035],seed[293],seed[3026],seed[973],seed[187],seed[364],seed[835],seed[1661],seed[3851],seed[3588],seed[3299],seed[3434],seed[4064],seed[3679],seed[2330],seed[1649],seed[3547],seed[829],seed[117],seed[2677],seed[1079],seed[890],seed[3999],seed[441],seed[3088],seed[4009],seed[2377],seed[1046],seed[2082],seed[1549],seed[3153],seed[1146],seed[2231],seed[240],seed[1754],seed[3274],seed[2912],seed[2532],seed[279],seed[1792],seed[3707],seed[1750],seed[853],seed[274],seed[2133],seed[3003],seed[1],seed[3624],seed[3879],seed[3281],seed[1404],seed[3615],seed[65],seed[2385],seed[4055],seed[327],seed[3595],seed[1173],seed[3568],seed[3766],seed[3917],seed[2378],seed[1242],seed[127],seed[1620],seed[248],seed[3076],seed[2370],seed[732],seed[768],seed[3012],seed[4020],seed[943],seed[391],seed[1346],seed[1968],seed[1100],seed[1912],seed[158],seed[2003],seed[963],seed[135],seed[3729],seed[2922],seed[306],seed[2886],seed[1807],seed[2100],seed[1533],seed[1347],seed[505],seed[108],seed[764],seed[543],seed[2814],seed[1487],seed[775],seed[982],seed[3496],seed[335],seed[1465],seed[1179],seed[3106],seed[1025],seed[3288],seed[1239],seed[150],seed[2490],seed[3930],seed[3481],seed[1475],seed[587],seed[2596],seed[499],seed[2919],seed[3951],seed[3259],seed[367],seed[3435],seed[1041],seed[3666],seed[2710],seed[2897],seed[1312],seed[2324],seed[1471],seed[235],seed[339],seed[736],seed[2862],seed[3969],seed[2264],seed[573],seed[1421],seed[1904],seed[1157],seed[3504],seed[2773],seed[1054],seed[1778],seed[3532],seed[358],seed[183],seed[2554],seed[159],seed[1826],seed[625],seed[1199],seed[1056],seed[2501],seed[2251],seed[1248],seed[2960],seed[233],seed[3285],seed[923],seed[453],seed[2277],seed[1731],seed[2030],seed[1640],seed[3018],seed[3296],seed[2907],seed[2848],seed[2858],seed[3114],seed[2625],seed[3245],seed[104],seed[983],seed[4015],seed[409],seed[173],seed[304],seed[2483],seed[3896],seed[1656],seed[1316],seed[3887],seed[3372],seed[3370],seed[3933],seed[2353],seed[1813],seed[3981],seed[3791],seed[2698],seed[2822],seed[374],seed[3864],seed[2332],seed[3498],seed[1823],seed[46],seed[1238],seed[1424],seed[3768],seed[3660],seed[2012],seed[1181],seed[1344],seed[354],seed[1696],seed[634],seed[1873],seed[1349],seed[604],seed[2614],seed[4095],seed[2772],seed[80],seed[3823],seed[3846],seed[3630],seed[1494],seed[1571],seed[2881],seed[3559],seed[3369],seed[947],seed[2079],seed[2801],seed[2013],seed[2075],seed[475],seed[2500],seed[351],seed[2362],seed[1410],seed[1155],seed[2693],seed[2418],seed[3730],seed[3636],seed[1270],seed[1204],seed[1838],seed[2191],seed[2867],seed[3137],seed[3847],seed[3811],seed[917],seed[1216],seed[699],seed[1379],seed[1715],seed[1215],seed[515],seed[1377],seed[1965],seed[3389],seed[1330],seed[1612],seed[578],seed[548],seed[3260],seed[3908],seed[3108],seed[3015],seed[1031],seed[1972],seed[517],seed[3099],seed[3415],seed[2080],seed[2600],seed[965],seed[1310],seed[3513],seed[1247],seed[2969],seed[1028],seed[2689],seed[880],seed[1191],seed[2093],seed[3125],seed[2830],seed[225],seed[3201],seed[3704],seed[3934],seed[16],seed[1634],seed[2208],seed[1752],seed[1858],seed[3665],seed[1140],seed[2847],seed[1060],seed[488],seed[2702],seed[1052],seed[856],seed[3071],seed[3198],seed[2258],seed[3512],seed[237],seed[2398],seed[785],seed[2589],seed[2416],seed[1250],seed[3393],seed[1417],seed[1072],seed[2587],seed[2544],seed[2853],seed[92],seed[1741],seed[495],seed[3954],seed[3265],seed[1489],seed[955],seed[1180],seed[1519],seed[1760],seed[1601],seed[1279],seed[522],seed[2563],seed[412],seed[2296],seed[772],seed[2197],seed[268],seed[996],seed[2417],seed[1177],seed[2891],seed[3312],seed[372],seed[2914],seed[3090],seed[2606],seed[597],seed[2234],seed[2743],seed[865],seed[1147],seed[1101],seed[3227],seed[4038],seed[3519],seed[2525],seed[203],seed[2005],seed[1524],seed[2738],seed[3255],seed[2269],seed[112],seed[378],seed[2709],seed[2413],seed[3204],seed[782],seed[3457],seed[2624],seed[3911],seed[1998],seed[1128],seed[1980],seed[4083],seed[4051],seed[2599],seed[1504],seed[1958],seed[139],seed[747],seed[3909],seed[945],seed[73],seed[3328],seed[3268],seed[1699],seed[2706],seed[2753],seed[2288],seed[2811],seed[3902],seed[353],seed[2887],seed[843],seed[629],seed[612],seed[2382],seed[371],seed[2036],seed[3349],seed[2827],seed[1009],seed[756],seed[2530],seed[1209],seed[418],seed[2303],seed[673],seed[152],seed[3667],seed[3622],seed[1567],seed[3244],seed[1672],seed[3362],seed[2227],seed[2989],seed[3680],seed[30],seed[1531],seed[2831],seed[2472],seed[3574],seed[496],seed[1911],seed[2463],seed[2641],seed[2846],seed[2312],seed[3617],seed[3813],seed[657],seed[1306],seed[3767],seed[1325],seed[2400],seed[1921],seed[2173],seed[821],seed[2562],seed[2216],seed[2719],seed[1774],seed[99],seed[3335],seed[21],seed[45],seed[3267],seed[1497],seed[2243],seed[678],seed[301],seed[2779],seed[177],seed[3266],seed[605],seed[1647],seed[2608],seed[1015],seed[2217],seed[129],seed[1971],seed[1881],seed[1722],seed[3145],seed[2894],seed[491],seed[868],seed[3477],seed[2177],seed[915],seed[3021],seed[2504],seed[3073],seed[3256],seed[1984],seed[1036],seed[163],seed[891],seed[1702],seed[106],seed[867],seed[2558],seed[161],seed[3154],seed[735],seed[1771],seed[419],seed[84],seed[1186],seed[3452],seed[3598],seed[2031],seed[1947],seed[3781],seed[3222],seed[993],seed[3403],seed[389],seed[2920],seed[2009],seed[3085],seed[1129],seed[3785],seed[136],seed[3777],seed[405],seed[3261],seed[125],seed[2311],seed[3809],seed[1010],seed[2864],seed[414],seed[803],seed[267],seed[3292],seed[4010],seed[426],seed[4001],seed[2308],seed[3190],seed[905],seed[3582],seed[2340],seed[916],seed[2615],seed[769],seed[3476],seed[1600],seed[3548],seed[1207],seed[784],seed[2179],seed[1548],seed[2749],seed[953],seed[75],seed[1520],seed[1986],seed[3807],seed[1227],seed[3377],seed[1530],seed[3619],seed[3871],seed[3678],seed[2223],seed[3893],seed[2358],seed[3338],seed[3282],seed[70],seed[3311],seed[197],seed[3765],seed[3497],seed[1832],seed[3763],seed[466],seed[1246],seed[3269],seed[3419],seed[3331],seed[3689],seed[2626],seed[4074],seed[1166],seed[3351],seed[714],seed[2091],seed[3200],seed[1755],seed[614],seed[1322],seed[3058],seed[3093],seed[198],seed[3038],seed[937],seed[1534],seed[3407],seed[833],seed[1910],seed[168],seed[2799],seed[2268],seed[4062],seed[1859],seed[1425],seed[3965],seed[2751],seed[3569],seed[2002],seed[705],seed[156],seed[3277],seed[3789],seed[2671],seed[1273],seed[2958],seed[3287],seed[1136],seed[3850],seed[470],seed[3516],seed[3994],seed[1159],seed[1780],seed[3884],seed[4086],seed[1788],seed[1418],seed[1735],seed[184],seed[3627],seed[1383],seed[2545],seed[2290],seed[2524],seed[2785],seed[540],seed[2705],seed[3501],seed[3410],seed[743],seed[1105],seed[2818],seed[751],seed[1450],seed[694],seed[385],seed[991],seed[1668],seed[3881],seed[3524],seed[2519],seed[3116],seed[1476],seed[3213],seed[2094],seed[2066],seed[1375],seed[3671],seed[2807],seed[901],seed[2637],seed[2437],seed[642],seed[3754],seed[2061],seed[2365],seed[428],seed[456],seed[4012],seed[1862],seed[3355],seed[1657],seed[1264],seed[3677],seed[911],seed[575],seed[1693],seed[2242],seed[3814],seed[1905],seed[1334],seed[3176],seed[3649],seed[1098],seed[878],seed[1937],seed[3308],seed[584],seed[455],seed[4017],seed[1506],seed[2513],seed[531],seed[1850],seed[67],seed[3946],seed[1773],seed[778],seed[2533],seed[3843],seed[3027],seed[3603],seed[2434],seed[1919],seed[3028],seed[660],seed[1670],seed[2065],seed[3511],seed[1111],seed[3531],seed[2499],seed[3128],seed[3517],seed[680],seed[1690],seed[2473],seed[2042],seed[4007],seed[284],seed[4054],seed[1700],seed[617],seed[381],seed[1522],seed[2457],seed[71],seed[704],seed[3290],seed[448],seed[2150],seed[3682],seed[2244],seed[3366],seed[1374],seed[4078],seed[2674],seed[3694],seed[733],seed[3885],seed[1762],seed[2298],seed[2849],seed[395],seed[3831],seed[930],seed[560],seed[3796],seed[1269],seed[145],seed[477],seed[2795],seed[3405],seed[3380],seed[3295],seed[794],seed[2798],seed[3998],seed[513],seed[1518],seed[877],seed[1062],seed[404],seed[1880],seed[1678],seed[3007],seed[3943],seed[3262],seed[1193],seed[3052],seed[2255],seed[1967],seed[1119],seed[3191],seed[2776],seed[554],seed[243],seed[1901],seed[783],seed[2343],seed[2364],seed[1305],seed[4046],seed[840],seed[2857],seed[3651],seed[3223],seed[606],seed[4079],seed[3988],seed[2595],seed[3749],seed[2474],seed[3949],seed[1370],seed[3054],seed[176],seed[1872],seed[3020],seed[3160],seed[2351],seed[2617],seed[645],seed[757],seed[1579],seed[2889],seed[2106],seed[2449],seed[717],seed[2609],seed[2583],seed[1688],seed[2520],seed[3805],seed[3985],seed[1350],seed[3102],seed[2904],seed[3983],seed[1134],seed[2316],seed[2739],seed[2412],seed[2445],seed[1295],seed[929],seed[651],seed[1358],seed[2976],seed[2636],seed[2399],seed[866],seed[3272],seed[1505],seed[3853],seed[2703],seed[121],seed[89],seed[1456],seed[1645],seed[3759],seed[2395],seed[1767],seed[386],seed[3728],seed[2837],seed[1890],seed[1074],seed[1663],seed[482],seed[1884],seed[2610],seed[3381],seed[689],seed[2593],seed[2730],seed[2431],seed[3738],seed[3004],seed[776],seed[3935],seed[640],seed[809],seed[557],seed[1263],seed[3105],seed[2538],seed[2429],seed[1113],seed[1145],seed[1491],seed[1420],seed[3558],seed[988],seed[656],seed[3066],seed[4053],seed[2004],seed[2816],seed[2843],seed[2982],seed[253],seed[47],seed[429],seed[2022],seed[2241],seed[1841],seed[2245],seed[1176],seed[3786],seed[3159],seed[2654],seed[2687],seed[2341],seed[4070],seed[2775],seed[3155],seed[402],seed[2833],seed[1684],seed[2376],seed[2212],seed[154],seed[2488],seed[2856],seed[708],seed[2446],seed[2371],seed[1103],seed[3898],seed[3238],seed[1787],seed[3747],seed[3829],seed[2804],seed[2096],seed[815],seed[261],seed[1732],seed[3037],seed[1390],seed[3376],seed[1856],seed[137],seed[60],seed[2784],seed[2211],seed[1597],seed[3748],seed[1055],seed[3621],seed[2224],seed[525],seed[532],seed[3987],seed[3462],seed[2270],seed[427],seed[3444],seed[479],seed[407],seed[2873],seed[3047],seed[147],seed[995],seed[669],seed[3359],seed[3095],seed[2424],seed[2306],seed[2660],seed[214],seed[2183],seed[181],seed[3952],seed[1964],seed[417],seed[2966],seed[2794],seed[828],seed[2971],seed[3620],seed[3314],seed[234],seed[3010],seed[486],seed[3554],seed[3278],seed[3711],seed[1818],seed[970],seed[2348],seed[1428],seed[3808],seed[969],seed[881],seed[4094],seed[3841],seed[1662],seed[897],seed[2238],seed[1564],seed[817],seed[4057],seed[2450],seed[1776],seed[3618],seed[3631],seed[2088],seed[3510],seed[1026],seed[1575],seed[4065],seed[72],seed[2696],seed[3801],seed[1568],seed[3566],seed[144],seed[3345],seed[2868],seed[1590],seed[2187],seed[4072],seed[478],seed[3608],seed[1626],seed[590],seed[41],seed[1449],seed[2359],seed[436],seed[442],seed[4089],seed[1630],seed[3192],seed[227],seed[2968],seed[2367],seed[3953],seed[1951],seed[1790],seed[3817],seed[1470],seed[4026],seed[3000],seed[56],seed[2152],seed[1139],seed[2451],seed[3334],seed[2931],seed[3367],seed[190],seed[847],seed[1464],seed[596],seed[862],seed[295],seed[3183],seed[17],seed[832],seed[3464],seed[1527],seed[1393],seed[872],seed[3703],seed[2077],seed[3827],seed[1577],seed[3408],seed[2250],seed[3576],seed[3305],seed[948],seed[773],seed[886],seed[1265],seed[1997],seed[2148],seed[1685],seed[4067],seed[3184],seed[1268],seed[1926],seed[2761],seed[1563],seed[3662],seed[2396],seed[3344],seed[1252],seed[2880],seed[437],seed[1466],seed[627],seed[762],seed[51],seed[842],seed[3293],seed[3068],seed[175],seed[839],seed[1763],seed[1051],seed[3894],seed[1460],seed[149],seed[2157],seed[469],seed[2550],seed[3440],seed[1949],seed[3420],seed[2384],seed[4037],seed[3873],seed[215],seed[1876],seed[2832],seed[357],seed[2374],seed[3571],seed[1090],seed[314],seed[2729],seed[2074],seed[4029],seed[3132],seed[3974],seed[1526],seed[912],seed[529],seed[2944],seed[1326],seed[1089],seed[3394],seed[1827],seed[3306],seed[3995],seed[413],seed[3616],seed[2305],seed[3836],seed[9],seed[4041],seed[1992],seed[1184],seed[3655],seed[2665],seed[1336],seed[2064],seed[3115],seed[81],seed[1586],seed[1272],seed[2200],seed[3418],seed[889],seed[3173],seed[1000],seed[3475],seed[1066],seed[2640],seed[503],seed[2825],seed[2192],seed[1073],seed[3856],seed[2139],seed[1885],seed[2040],seed[254],seed[2821],seed[2167],seed[547],seed[1032],seed[3575],seed[591],seed[2136],seed[1226],seed[3962],seed[1908],seed[471],seed[4068],seed[3357],seed[2205],seed[282],seed[3368],seed[3432],seed[3469],seed[272],seed[2226],seed[180],seed[3990],seed[1160],seed[1037],seed[2062],seed[1679],seed[487],seed[3092],seed[2199],seed[3083],seed[1473],seed[1742],seed[2476],seed[820],seed[1122],seed[3762],seed[217],seed[375],seed[2796],seed[4033],seed[2198],seed[1582],seed[1212],seed[3800],seed[2168],seed[3196],seed[162],seed[2056],seed[1245],seed[2310],seed[4],seed[2259],seed[3866],seed[2309],seed[1389],seed[3329],seed[2302],seed[2470],seed[3997],seed[2497],seed[2789],seed[2731],seed[2611],seed[1003],seed[4022],seed[3426],seed[160],seed[2783],seed[23],seed[2733],seed[1913],seed[3538],seed[2990],seed[3117],seed[3107],seed[537],seed[2381],seed[3710],seed[2453],seed[1502],seed[1723],seed[1384],seed[1772],seed[1902],seed[3333],seed[985],seed[3110],seed[3604],seed[1673],seed[3597],seed[2656],seed[1743],seed[20],seed[1353],seed[1485],seed[3216],seed[1785],seed[3316],seed[1366],seed[693],seed[3546],seed[3875],seed[1102],seed[2882],seed[4011],seed[3019],seed[3986],seed[3633],seed[1260],seed[1831],seed[706],seed[3103],seed[2254],seed[3398],seed[3025],seed[526],seed[3141],seed[3024],seed[3977],seed[2566],seed[3307],seed[1220],seed[826],seed[323],seed[1583],seed[3727],seed[2182],seed[810],seed[1650],seed[224],seed[1321],seed[2142],seed[283],seed[2054],seed[3294],seed[2741],seed[2620],seed[1092],seed[2027],seed[2716],seed[1369],seed[483],seed[715],seed[7],seed[2915],seed[3143],seed[2007],seed[3482],seed[1455],seed[2515],seed[2475],seed[126],seed[990],seed[91],seed[103],seed[992],seed[2176],seed[1532],seed[2045],seed[2456],seed[586],seed[1618],seed[3925],seed[932],seed[3761],seed[3313],seed[1376],seed[1692],seed[3354],seed[2404],seed[1596],seed[755],seed[3382],seed[709],seed[687],seed[2537],seed[3506],seed[2252],seed[2844],seed[1570],seed[580],seed[2746],seed[2117],seed[2145],seed[2684],seed[50],seed[888],seed[100],seed[3422],seed[3343],seed[887],seed[1955],seed[1782],seed[2954],seed[3241],seed[2059],seed[2084],seed[2166],seed[3330],seed[787],seed[3882],seed[3507],seed[1462],seed[1695],seed[523],seed[3553],seed[1192],seed[2999],seed[3412],seed[1415],seed[3219],seed[1423],seed[4056],seed[1099],seed[3876],seed[1283],seed[1198],seed[324],seed[2754],seed[3672],seed[3741],seed[1639],seed[677],seed[1256],seed[3158],seed[2855],seed[3659],seed[770],seed[4063],seed[3171],seed[962],seed[232],seed[2228],seed[1371],seed[55],seed[1029],seed[1234],seed[3541],seed[1698],seed[3119],seed[1886],seed[3347],seed[1629],seed[1825],seed[4082],seed[1615],seed[2337],seed[281],seed[507],seed[3858],seed[570],seed[128],seed[271],seed[1953],seed[3611],seed[430],seed[3522],seed[2560],seed[2745],seed[2097],seed[3750],seed[519],seed[3653],seed[1258],seed[1278],seed[3534],seed[1472],seed[1352],seed[1703],seed[2720],seed[1830],seed[2246],seed[2435],seed[3956],seed[3932],seed[1075],seed[510],seed[216],seed[2350],seed[2235],seed[545],seed[4040],seed[2762],seed[255],seed[3414],seed[1554],seed[2974],seed[276],seed[1900],seed[490],seed[392]}),
        .cross_prob(cross_prob),
        .codeword(codeword3),
        .received(received3)
        );
    
    bsc bsc4(
        .clk(clk),
        .reset(reset),
        .seed({seed[3009],seed[3046],seed[268],seed[200],seed[1455],seed[1031],seed[3307],seed[3096],seed[3119],seed[493],seed[2671],seed[1150],seed[3621],seed[412],seed[3785],seed[2453],seed[2034],seed[3350],seed[3498],seed[3598],seed[2570],seed[3979],seed[1970],seed[902],seed[847],seed[791],seed[1309],seed[404],seed[130],seed[3735],seed[39],seed[1737],seed[3400],seed[3817],seed[3111],seed[2839],seed[3921],seed[3813],seed[3623],seed[1674],seed[3746],seed[4073],seed[483],seed[3831],seed[1110],seed[1806],seed[1384],seed[429],seed[1207],seed[1091],seed[960],seed[749],seed[2389],seed[1360],seed[3195],seed[3468],seed[3728],seed[3044],seed[713],seed[1498],seed[1263],seed[155],seed[3033],seed[3857],seed[3691],seed[1247],seed[1220],seed[2747],seed[3557],seed[1715],seed[562],seed[7],seed[3408],seed[1506],seed[3646],seed[2065],seed[2864],seed[2422],seed[1611],seed[3045],seed[4093],seed[1854],seed[1914],seed[2167],seed[2125],seed[1616],seed[2481],seed[2889],seed[569],seed[4080],seed[2812],seed[987],seed[549],seed[2134],seed[1516],seed[1284],seed[2782],seed[3030],seed[2693],seed[278],seed[1158],seed[3308],seed[3690],seed[3438],seed[3624],seed[2666],seed[2713],seed[1833],seed[1820],seed[2676],seed[12],seed[1633],seed[2658],seed[335],seed[542],seed[2925],seed[1470],seed[3609],seed[574],seed[3645],seed[3605],seed[2896],seed[3680],seed[2630],seed[2610],seed[897],seed[3227],seed[3364],seed[2221],seed[2386],seed[3975],seed[903],seed[2979],seed[3015],seed[3633],seed[3058],seed[2201],seed[399],seed[1156],seed[2659],seed[1035],seed[3446],seed[1074],seed[820],seed[193],seed[3882],seed[3516],seed[3991],seed[1818],seed[2541],seed[2060],seed[666],seed[2727],seed[71],seed[660],seed[3504],seed[3913],seed[99],seed[3283],seed[2072],seed[3812],seed[3767],seed[3532],seed[3346],seed[1234],seed[1959],seed[450],seed[3077],seed[14],seed[1505],seed[3614],seed[1204],seed[817],seed[1072],seed[1011],seed[1965],seed[596],seed[3951],seed[1051],seed[2147],seed[174],seed[2656],seed[804],seed[2959],seed[3215],seed[98],seed[1194],seed[3117],seed[1332],seed[2490],seed[3715],seed[2780],seed[2950],seed[2878],seed[3640],seed[1856],seed[708],seed[3788],seed[3322],seed[2370],seed[1657],seed[1655],seed[838],seed[2249],seed[423],seed[1721],seed[2188],seed[2772],seed[2967],seed[1105],seed[869],seed[3319],seed[2771],seed[4016],seed[2619],seed[711],seed[1858],seed[3896],seed[3368],seed[1756],seed[242],seed[3945],seed[2206],seed[2230],seed[572],seed[3681],seed[2280],seed[181],seed[2284],seed[1160],seed[116],seed[2058],seed[3189],seed[3796],seed[2894],seed[637],seed[754],seed[1282],seed[742],seed[1040],seed[766],seed[1980],seed[2668],seed[2421],seed[3310],seed[2269],seed[59],seed[182],seed[2555],seed[165],seed[682],seed[1705],seed[2022],seed[1998],seed[491],seed[400],seed[720],seed[3964],seed[2568],seed[3130],seed[2567],seed[2688],seed[2363],seed[1610],seed[1813],seed[1411],seed[2311],seed[2182],seed[3049],seed[1169],seed[3328],seed[3843],seed[3141],seed[1971],seed[1672],seed[306],seed[2024],seed[2351],seed[1266],seed[3860],seed[1739],seed[2665],seed[3198],seed[1500],seed[3657],seed[2867],seed[3747],seed[2973],seed[1094],seed[3769],seed[566],seed[1413],seed[2775],seed[2640],seed[3494],seed[3205],seed[1932],seed[3097],seed[593],seed[3886],seed[3524],seed[2598],seed[1210],seed[1696],seed[2604],seed[3210],seed[3039],seed[492],seed[2863],seed[60],seed[1188],seed[1767],seed[1319],seed[3406],seed[3658],seed[4090],seed[2834],seed[2457],seed[1477],seed[2859],seed[272],seed[1046],seed[3148],seed[2492],seed[4060],seed[2231],seed[934],seed[203],seed[1133],seed[2124],seed[967],seed[4046],seed[386],seed[294],seed[2911],seed[845],seed[169],seed[2448],seed[1253],seed[2919],seed[3707],seed[3465],seed[223],seed[1771],seed[1568],seed[3556],seed[2339],seed[1810],seed[1629],seed[2736],seed[420],seed[3334],seed[1566],seed[2843],seed[1837],seed[2399],seed[3485],seed[19],seed[786],seed[3798],seed[725],seed[1957],seed[3125],seed[102],seed[2813],seed[931],seed[3804],seed[1244],seed[1028],seed[3694],seed[1059],seed[3577],seed[1060],seed[2025],seed[119],seed[1324],seed[1826],seed[1708],seed[2765],seed[2857],seed[3288],seed[570],seed[737],seed[1951],seed[2452],seed[3380],seed[1750],seed[3123],seed[115],seed[787],seed[662],seed[2160],seed[878],seed[834],seed[1054],seed[2810],seed[531],seed[1396],seed[263],seed[3133],seed[82],seed[1488],seed[3825],seed[2478],seed[113],seed[597],seed[507],seed[2085],seed[1277],seed[3171],seed[2877],seed[108],seed[2573],seed[776],seed[1988],seed[703],seed[3875],seed[994],seed[2648],seed[2028],seed[2184],seed[3375],seed[527],seed[3251],seed[3729],seed[1982],seed[3292],seed[2396],seed[151],seed[3844],seed[3655],seed[137],seed[3669],seed[1180],seed[627],seed[2788],seed[1582],seed[2687],seed[138],seed[2113],seed[1978],seed[2050],seed[2094],seed[187],seed[1387],seed[831],seed[40],seed[316],seed[1489],seed[3683],seed[3572],seed[112],seed[2618],seed[854],seed[4044],seed[460],seed[1814],seed[362],seed[500],seed[3930],seed[2700],seed[2714],seed[3803],seed[1595],seed[1435],seed[215],seed[2794],seed[1975],seed[674],seed[2491],seed[1699],seed[3137],seed[1613],seed[3032],seed[3037],seed[2070],seed[3706],seed[3667],seed[3642],seed[1353],seed[135],seed[2271],seed[332],seed[2985],seed[1355],seed[1403],seed[1995],seed[396],seed[3026],seed[2746],seed[219],seed[2236],seed[2251],seed[3947],seed[794],seed[1122],seed[31],seed[3588],seed[1786],seed[3933],seed[3379],seed[3267],seed[675],seed[41],seed[3443],seed[1599],seed[545],seed[2850],seed[3279],seed[1717],seed[3779],seed[52],seed[2807],seed[1539],seed[3997],seed[3617],seed[1231],seed[2735],seed[914],seed[1996],seed[3344],seed[3],seed[1223],seed[986],seed[702],seed[2402],seed[663],seed[563],seed[205],seed[1893],seed[2703],seed[2970],seed[671],seed[2243],seed[454],seed[1077],seed[2498],seed[2130],seed[1392],seed[1926],seed[74],seed[1409],seed[1546],seed[3156],seed[3473],seed[1412],seed[3873],seed[1337],seed[3404],seed[3878],seed[1747],seed[1943],seed[3418],seed[2063],seed[315],seed[1710],seed[23],seed[1183],seed[2319],seed[3464],seed[2942],seed[760],seed[4010],seed[2729],seed[2082],seed[1394],seed[941],seed[2428],seed[1153],seed[2384],seed[1646],seed[2446],seed[378],seed[3794],seed[1000],seed[1440],seed[3135],seed[3491],seed[3518],seed[3188],seed[3241],seed[1395],seed[1671],seed[3839],seed[2616],seed[3471],seed[2226],seed[2318],seed[3434],seed[3374],seed[2196],seed[325],seed[3560],seed[1637],seed[937],seed[1200],seed[1476],seed[946],seed[285],seed[2220],seed[2677],seed[624],seed[3367],seed[431],seed[3534],seed[3291],seed[3385],seed[3566],seed[3676],seed[1424],seed[1844],seed[3682],seed[3100],seed[2008],seed[3178],seed[598],seed[107],seed[1534],seed[2509],seed[1731],seed[3483],seed[3738],seed[1380],seed[2081],seed[1149],seed[1103],seed[199],seed[2029],seed[2769],seed[1299],seed[2732],seed[3259],seed[1132],seed[406],seed[3474],seed[1625],seed[1684],seed[3318],seed[976],seed[3731],seed[3153],seed[1903],seed[626],seed[2617],seed[188],seed[680],seed[2635],seed[331],seed[640],seed[829],seed[3463],seed[526],seed[401],seed[2720],seed[3104],seed[2503],seed[1556],seed[1925],seed[3508],seed[1704],seed[437],seed[3819],seed[2836],seed[347],seed[1827],seed[373],seed[345],seed[3601],seed[1983],seed[3360],seed[3711],seed[4089],seed[1084],seed[1316],seed[288],seed[3127],seed[938],seed[573],seed[2062],seed[28],seed[3495],seed[3923],seed[1920],seed[1614],seed[581],seed[2380],seed[1467],seed[745],seed[1656],seed[3401],seed[1673],seed[571],seed[2208],seed[3759],seed[2451],seed[3266],seed[1290],seed[1789],seed[1669],seed[217],seed[1512],seed[2036],seed[2071],seed[1269],seed[1843],seed[51],seed[2104],seed[2033],seed[1991],seed[2506],seed[3685],seed[1466],seed[1388],seed[4088],seed[1815],seed[1691],seed[2578],seed[706],seed[3582],seed[2204],seed[3229],seed[1085],seed[432],seed[2832],seed[3220],seed[3000],seed[1437],seed[158],seed[2296],seed[2507],seed[621],seed[3751],seed[171],seed[2173],seed[2300],seed[3031],seed[2107],seed[2288],seed[1964],seed[2642],seed[1563],seed[1897],seed[1499],seed[783],seed[3602],seed[3632],seed[1314],seed[3353],seed[18],seed[3616],seed[2809],seed[314],seed[3919],seed[1758],seed[3703],seed[3708],seed[2193],seed[1538],seed[2789],seed[1801],seed[4082],seed[2073],seed[2279],seed[1921],seed[81],seed[2026],seed[1723],seed[1013],seed[1587],seed[3166],seed[2934],seed[865],seed[1361],seed[2995],seed[653],seed[2006],seed[2390],seed[1834],seed[3073],seed[899],seed[2234],seed[2624],seed[966],seed[407],seed[2157],seed[66],seed[2023],seed[812],seed[3580],seed[300],seed[380],seed[1985],seed[1639],seed[3720],seed[3845],seed[1586],seed[4064],seed[2368],seed[1227],seed[3496],seed[4071],seed[3705],seed[2653],seed[3349],seed[2487],seed[3074],seed[3576],seed[3355],seed[456],seed[2767],seed[3841],seed[2808],seed[411],seed[1630],seed[616],seed[1064],seed[13],seed[2414],seed[2566],seed[1167],seed[3814],seed[1778],seed[2672],seed[1911],seed[633],seed[9],seed[1176],seed[1181],seed[1930],seed[991],seed[2704],seed[832],seed[3523],seed[2643],seed[3078],seed[1864],seed[1529],seed[3853],seed[1113],seed[2981],seed[2999],seed[2890],seed[789],seed[2185],seed[179],seed[1260],seed[3174],seed[942],seed[1255],seed[2098],seed[2538],seed[1447],seed[308],seed[1627],seed[1137],seed[270],seed[1553],seed[3143],seed[185],seed[3414],seed[2644],seed[3154],seed[2429],seed[2454],seed[814],seed[3028],seed[3884],seed[1984],seed[2365],seed[1608],seed[1565],seed[1313],seed[910],seed[874],seed[2350],seed[3020],seed[591],seed[1386],seed[3990],seed[416],seed[1206],seed[2357],seed[1677],seed[1949],seed[3625],seed[291],seed[2702],seed[2623],seed[1326],seed[45],seed[344],seed[2483],seed[1584],seed[2929],seed[3219],seed[361],seed[3088],seed[2077],seed[235],seed[430],seed[1675],seed[2021],seed[1762],seed[1787],seed[3543],seed[1693],seed[2560],seed[3584],seed[3282],seed[844],seed[143],seed[3050],seed[307],seed[3341],seed[1146],seed[42],seed[3943],seed[1760],seed[2632],seed[3208],seed[3330],seed[722],seed[3949],seed[2508],seed[402],seed[1759],seed[1436],seed[2348],seed[4053],seed[2444],seed[922],seed[908],seed[3458],seed[1378],seed[3663],seed[1623],seed[871],seed[3196],seed[1768],seed[3252],seed[305],seed[3451],seed[3752],seed[1752],seed[2575],seed[2800],seed[1010],seed[3072],seed[2387],seed[2546],seed[1919],seed[2158],seed[718],seed[679],seed[3757],seed[2440],seed[4050],seed[227],seed[3835],seed[781],seed[1119],seed[2456],seed[2980],seed[3678],seed[3739],seed[2937],seed[2759],seed[1907],seed[3548],seed[474],seed[3336],seed[1992],seed[583],seed[1179],seed[3679],seed[417],seed[1860],seed[4079],seed[2493],seed[1873],seed[2106],seed[2138],seed[3014],seed[2516],seed[2057],seed[3022],seed[1067],seed[1532],seed[1274],seed[588],seed[3129],seed[2791],seed[3865],seed[122],seed[1092],seed[1017],seed[2891],seed[3164],seed[958],seed[2885],seed[2069],seed[1257],seed[1915],seed[1159],seed[4014],seed[1305],seed[3562],seed[1716],seed[2627],seed[2056],seed[2340],seed[2172],seed[148],seed[3057],seed[3297],seed[2922],seed[2292],seed[3957],seed[97],seed[128],seed[2753],seed[3052],seed[3412],seed[2673],seed[3920],seed[575],seed[201],seed[1665],seed[520],seed[3699],seed[1405],seed[2913],seed[2792],seed[77],seed[3388],seed[395],seed[2406],seed[144],seed[4028],seed[2531],seed[3828],seed[2449],seed[3898],seed[2411],seed[4055],seed[3615],seed[2636],seed[1558],seed[560],seed[2347],seed[2683],seed[1340],seed[133],seed[2797],seed[732],seed[2997],seed[2593],seed[2317],seed[819],seed[2301],seed[296],seed[3488],seed[1829],seed[3982],seed[2730],seed[3124],seed[534],seed[2032],seed[763],seed[816],seed[1668],seed[1927],seed[2222],seed[1901],seed[3537],seed[3575],seed[1761],seed[289],seed[3186],seed[2198],seed[222],seed[1371],seed[2825],seed[601],seed[777],seed[2191],seed[3940],seed[2875],seed[2265],seed[1987],seed[3815],seed[3163],seed[391],seed[3559],seed[2978],seed[4],seed[2447],seed[72],seed[2123],seed[3637],seed[95],seed[1681],seed[1811],seed[3758],seed[2048],seed[240],seed[3594],seed[2295],seed[2831],seed[2581],seed[3043],seed[2410],seed[3824],seed[2007],seed[1006],seed[1724],seed[2953],seed[2404],seed[3054],seed[1809],seed[2849],seed[343],seed[1358],seed[1288],seed[3326],seed[4002],seed[2290],seed[1391],seed[1254],seed[940],seed[25],seed[2725],seed[644],seed[2115],seed[3021],seed[4067],seed[1297],seed[372],seed[2341],seed[1635],seed[3644],seed[3478],seed[1294],seed[3607],seed[4052],seed[2315],seed[1147],seed[350],seed[4026],seed[3149],seed[2038],seed[2031],seed[780],seed[697],seed[2822],seed[1869],seed[1221],seed[3320],seed[3958],seed[1766],seed[1184],seed[1136],seed[1644],seed[3626],seed[1486],seed[1754],seed[2096],seed[1302],seed[1480],seed[4017],seed[4035],seed[3927],seed[1116],seed[916],seed[1770],seed[2707],seed[1536],seed[1036],seed[3253],seed[1963],seed[3880],seed[2272],seed[3999],seed[1757],seed[2872],seed[694],seed[4062],seed[2554],seed[1725],seed[3959],seed[2010],seed[1073],seed[988],seed[252],seed[2586],seed[3695],seed[3363],seed[2824],seed[1709],seed[1414],seed[2544],seed[3545],seed[1654],seed[1946],seed[3142],seed[1020],seed[1393],seed[1454],seed[2542],seed[1289],seed[2256],seed[959],seed[1268],seed[304],seed[759],seed[79],seed[3549],seed[2382],seed[2883],seed[4038],seed[3387],seed[2171],seed[3005],seed[3883],seed[2267],seed[3087],seed[2726],seed[1124],seed[3976],seed[1853],seed[709],seed[1792],seed[1069],seed[211],seed[3442],seed[3937],seed[2018],seed[394],seed[3131],seed[1492],seed[896],seed[849],seed[214],seed[2868],seed[1323],seed[2461],seed[951],seed[2691],seed[3296],seed[3567],seed[3204],seed[815],seed[1056],seed[3306],seed[1632],seed[62],seed[1478],seed[2227],seed[3822],seed[3132],seed[3324],seed[172],seed[3102],seed[3082],seed[1940],seed[756],seed[194],seed[2881],seed[2907],seed[850],seed[2355],seed[1518],seed[249],seed[2670],seed[3247],seed[837],seed[2304],seed[843],seed[1218],seed[1249],seed[2572],seed[359],seed[3106],seed[3277],seed[2738],seed[298],seed[618],seed[2177],seed[2611],seed[3152],seed[2327],seed[856],seed[3255],seed[1857],seed[3583],seed[2470],seed[700],seed[2874],seed[579],seed[1631],seed[1032],seed[1166],seed[3926],seed[3370],seed[3709],seed[2294],seed[397],seed[836],seed[3238],seed[351],seed[3954],seed[2988],seed[1193],seed[1842],seed[1406],seed[3784],seed[3972],seed[2019],seed[2882],seed[1390],seed[1485],seed[1344],seed[2450],seed[2179],seed[2706],seed[1592],seed[2579],seed[2401],seed[2674],seed[2424],seed[311],seed[891],seed[1976],seed[2375],seed[2865],seed[2485],seed[1428],seed[3659],seed[1471],seed[1561],seed[2212],seed[3864],seed[355],seed[3352],seed[2900],seed[3486],seed[446],seed[1776],seed[1177],seed[568],seed[2861],seed[488],seed[2061],seed[2281],seed[465],seed[2165],seed[654],seed[2606],seed[2285],seed[1140],seed[2298],seed[1900],seed[3335],seed[3967],seed[911],seed[731],seed[2910],seed[164],seed[348],seed[2047],seed[1451],seed[1549],seed[1560],seed[912],seed[150],seed[3953],seed[312],seed[225],seed[243],seed[3487],seed[999],seed[953],seed[1504],seed[747],seed[730],seed[497],seed[1415],seed[3236],seed[3298],seed[1507],seed[2142],seed[3956],seed[2701],seed[75],seed[1062],seed[485],seed[1401],seed[1846],seed[2187],seed[2960],seed[3774],seed[3396],seed[673],seed[717],seed[1431],seed[1003],seed[3382],seed[1913],seed[3521],seed[580],seed[1527],seed[2975],seed[1267],seed[2535],seed[3966],seed[2828],seed[1198],seed[3517],seed[3889],seed[3454],seed[2425],seed[522],seed[161],seed[933],seed[3772],seed[1604],seed[1692],seed[1154],seed[876],seed[3730],seed[3475],seed[2639],seed[641],seed[1531],seed[2823],seed[811],seed[3365],seed[2846],seed[2525],seed[512],seed[3847],seed[3497],seed[3526],seed[1502],seed[2645],seed[585],seed[2592],seed[398],seed[1535],seed[525],seed[3193],seed[603],seed[1670],seed[2122],seed[3392],seed[3946],seed[24],seed[1107],seed[3998],seed[2916],seed[1058],seed[35],seed[748],seed[1803],seed[1589],seed[2600],seed[2977],seed[2009],seed[1548],seed[4015],seed[36],seed[1667],seed[3762],seed[2228],seed[436],seed[2091],seed[689],seed[2126],seed[3460],seed[2499],seed[3608],seed[2376],seed[1005],seed[4083],seed[3978],seed[4030],seed[3915],seed[3677],seed[2553],seed[3323],seed[2286],seed[89],seed[605],seed[1063],seed[1261],seed[2150],seed[1783],seed[1134],seed[2949],seed[602],seed[521],seed[746],seed[3697],seed[1640],seed[3151],seed[2426],seed[3359],seed[1443],seed[247],seed[2246],seed[2373],seed[620],seed[632],seed[455],seed[1609],seed[1322],seed[3611],seed[1519],seed[392],seed[1039],seed[3931],seed[121],seed[617],seed[2833],seed[1753],seed[145],seed[1205],seed[197],seed[2011],seed[1278],seed[1408],seed[178],seed[977],seed[1938],seed[2076],seed[2276],seed[3118],seed[3212],seed[2930],seed[3634],seed[2921],seed[638],seed[1571],seed[297],seed[2099],seed[2948],seed[3013],seed[3453],seed[949],seed[443],seed[2169],seed[303],seed[1969],seed[2958],seed[3895],seed[2408],seed[1429],seed[2001],seed[232],seed[1937],seed[2998],seed[2563],seed[807],seed[1475],seed[1482],seed[3639],seed[1400],seed[2596],seed[2705],seed[890],seed[375],seed[3808],seed[2915],seed[1374],seed[1840],seed[1318],seed[3996],seed[3126],seed[882],seed[950],seed[2074],seed[1093],seed[1583],seed[3300],seed[4074],seed[3613],seed[924],seed[1962],seed[2328],seed[965],seed[3520],seed[3619],seed[3529],seed[2143],seed[3175],seed[1680],seed[228],seed[466],seed[508],seed[2080],seed[2313],seed[2200],seed[650],seed[1125],seed[2356],seed[3936],seed[4004],seed[1083],seed[858],seed[1349],seed[3373],seed[1698],seed[209],seed[3698],seed[3971],seed[1389],seed[2003],seed[3903],seed[1043],seed[3109],seed[3989],seed[2893],seed[2040],seed[2244],seed[505],seed[2178],seed[576],seed[353],seed[3285],seed[2764],seed[91],seed[1356],seed[1808],seed[3112],seed[2161],seed[3480],seed[728],seed[607],seed[4066],seed[1430],seed[3832],seed[3554],seed[1816],seed[2545],seed[652],seed[1828],seed[271],seed[2240],seed[3047],seed[274],seed[3017],seed[2936],seed[1121],seed[877],seed[2684],seed[346],seed[2128],seed[2964],seed[1434],seed[1694],seed[87],seed[424],seed[1591],seed[3356],seed[114],seed[822],seed[1262],seed[2982],seed[1600],seed[2164],seed[3809],seed[4006],seed[1233],seed[3856],seed[913],seed[3775],seed[2361],seed[2739],seed[1372],seed[467],seed[770],seed[1450],seed[2109],seed[3603],seed[661],seed[2966],seed[3377],seed[2250],seed[4047],seed[655],seed[608],seed[1222],seed[969],seed[2842],seed[3648],seed[494],seed[239],seed[909],seed[2030],seed[687],seed[3091],seed[1848],seed[3618],seed[2901],seed[32],seed[715],seed[496],seed[166],seed[926],seed[1228],seed[1805],seed[4091],seed[2420],seed[3984],seed[1933],seed[901],seed[139],seed[830],seed[2749],seed[2170],seed[3098],seed[3718],seed[2695],seed[3362],seed[2622],seed[2441],seed[769],seed[469],seed[2145],seed[2235],seed[801],seed[1474],seed[1928],seed[2879],seed[1765],seed[3421],seed[1178],seed[1835],seed[1420],seed[3834],seed[2612],seed[1590],seed[3675],seed[2757],seed[1606],seed[3952],seed[3278],seed[755],seed[3941],seed[84],seed[1774],seed[963],seed[2273],seed[2131],seed[900],seed[1296],seed[2078],seed[3852],seed[905],seed[1238],seed[1989],seed[2652],seed[1624],seed[1009],seed[2105],seed[490],seed[3234],seed[1023],seed[2924],seed[1544],seed[1034],seed[4007],seed[936],seed[3547],seed[561],seed[3327],seed[3668],seed[1375],seed[4018],seed[69],seed[3888],seed[2268],seed[1952],seed[3505],seed[2391],seed[883],seed[1312],seed[3386],seed[3674],seed[2364],seed[613],seed[471],seed[1866],seed[2946],seed[1095],seed[2751],seed[3622],seed[1821],seed[555],seed[2895],seed[3851],seed[1917],seed[978],seed[1243],seed[805],seed[1330],seed[2067],seed[1979],seed[3961],seed[1345],seed[2603],seed[3411],seed[2637],seed[1799],seed[3413],seed[4000],seed[3258],seed[886],seed[2093],seed[157],seed[1219],seed[948],seed[1252],seed[3546],seed[3665],seed[3743],seed[3929],seed[3912],seed[3908],seed[584],seed[586],seed[125],seed[1785],seed[3140],seed[1459],seed[3760],seed[1742],seed[1626],seed[3745],seed[1923],seed[3089],seed[442],seed[2349],seed[67],seed[2087],seed[3254],seed[2302],seed[1797],seed[2345],seed[3136],seed[1075],seed[1327],seed[1540],seed[635],seed[2761],seed[3818],seed[1550],seed[3450],seed[881],seed[3407],seed[253],seed[1720],seed[2504],seed[3110],seed[301],seed[1385],seed[363],seed[1891],seed[2909],seed[317],seed[547],seed[511],seed[639],seed[2935],seed[3604],seed[1916],seed[2316],seed[1029],seed[3426],seed[772],seed[1446],seed[2260],seed[2321],seed[594],seed[326],seed[3983],seed[3565],seed[3733],seed[729],seed[3850],seed[2785],seed[3969],seed[3416],seed[664],seed[3347],seed[1612],seed[688],seed[2466],seed[3391],seed[3977],seed[3939],seed[3811],seed[1007],seed[3686],seed[379],seed[2016],seed[3980],seed[2951],seed[3402],seed[928],seed[3489],seed[322],seed[2431],seed[767],seed[2395],seed[230],seed[1303],seed[3748],seed[3906],seed[921],seed[221],seed[3661],seed[510],seed[1666],seed[1473],seed[3008],seed[1650],seed[3061],seed[147],seed[3466],seed[458],seed[3372],seed[686],seed[1906],seed[3872],seed[1264],seed[1120],seed[384],seed[3243],seed[2569],seed[1687],seed[866],seed[556],seed[2477],seed[724],seed[980],seed[2550],seed[409],seed[917],seed[3771],seed[1555],seed[2608],seed[1185],seed[589],seed[3034],seed[216],seed[2468],seed[2657],seed[647],seed[2803],seed[1643],seed[2059],seed[2101],seed[1298],seed[2042],seed[3176],seed[3993],seed[1364],seed[971],seed[3717],seed[1607],seed[68],seed[2781],seed[2920],seed[1245],seed[1711],seed[1562],seed[3654],seed[1494],seed[3287],seed[282],seed[1187],seed[1730],seed[309],seed[2561],seed[2799],seed[3786],seed[1577],seed[2841],seed[699],seed[1905],seed[2638],seed[4095],seed[3509],seed[1781],seed[2559],seed[2602],seed[149],seed[117],seed[1004],seed[3740],seed[3535],seed[2941],seed[1367],seed[1572],seed[788],seed[1291],seed[1664],seed[302],seed[930],seed[207],seed[751],seed[1130],seed[719],seed[2479],seed[3606],seed[1888],seed[3250],seed[1745],seed[2181],seed[1129],seed[3085],seed[275],seed[2218],seed[735],seed[1131],seed[2917],seed[3261],seed[4022],seed[390],seed[1918],seed[1163],seed[109],seed[448],seed[3826],seed[2151],seed[2027],seed[90],seed[3536],seed[2938],seed[1143],seed[3122],seed[377],seed[543],seed[495],seed[1079],seed[3628],seed[472],seed[177],seed[1071],seed[3684],seed[3120],seed[1875],seed[1172],seed[3514],seed[3165],seed[2084],seed[875],seed[3948],seed[3286],seed[3573],seed[4057],seed[356],seed[4019],seed[3909],seed[504],seed[3827],seed[1295],seed[57],seed[860],seed[3419],seed[3209],seed[2360],seed[3029],seed[3477],seed[4008],seed[1567],seed[170],seed[3002],seed[2342],seed[2562],seed[58],seed[1662],seed[3482],seed[2811],seed[984],seed[3519],seed[3224],seed[2472],seed[393],seed[428],seed[3035],seed[3256],seed[2183],seed[2203],seed[2053],seed[2320],seed[3274],seed[611],seed[658],seed[2523],seed[710],seed[1645],seed[2412],seed[3312],seed[3228],seed[2745],seed[1369],seed[1794],seed[281],seed[2871],seed[1986],seed[3018],seed[2821],seed[1545],seed[774],seed[4020],seed[3260],seed[636],seed[1037],seed[1763],seed[2192],seed[907],seed[2862],seed[544],seed[761],seed[2718],seed[1239],seed[1022],seed[4045],seed[2679],seed[2983],seed[1523],seed[2002],seed[3108],seed[3447],seed[3113],seed[3636],seed[3599],seed[993],seed[1108],seed[3870],seed[123],seed[2787],seed[3430],seed[167],seed[1735],seed[532],seed[3290],seed[3492],seed[146],seed[683],seed[892],seed[2486],seed[919],seed[685],seed[2912],seed[2888],seed[3742],seed[1270],seed[1772],seed[2464],seed[3284],seed[990],seed[2796],seed[1283],seed[1881],seed[1990],seed[2004],seed[389],seed[1524],seed[105],seed[1216],seed[1647],seed[853],seed[3476],seed[2136],seed[1511],seed[3202],seed[1841],seed[1484],seed[1383],seed[3107],seed[813],seed[1559],seed[3265],seed[435],seed[3099],seed[3422],seed[2918],seed[1338],seed[295],seed[1379],seed[3144],seed[524],seed[3805],seed[2664],seed[1968],seed[3182],seed[2969],seed[1065],seed[2584],seed[2580],seed[3056],seed[1462],seed[894],seed[1936],seed[3836],seed[1569],seed[2309],seed[1086],seed[3019],seed[4025],seed[425],seed[3833],seed[2906],seed[365],seed[2991],seed[3539],seed[1135],seed[2518],seed[1885],seed[1743],seed[1839],seed[2369],seed[864],seed[2520],seed[3242],seed[1448],seed[56],seed[333],seed[4043],seed[76],seed[83],seed[1780],seed[352],seed[3838],seed[2416],seed[369],seed[1317],seed[1142],seed[2766],seed[3462],seed[806],seed[2529],seed[3369],seed[37],seed[3907],seed[2536],seed[3868],seed[590],seed[2710],seed[2495],seed[1495],seed[2140],seed[2721],seed[3249],seed[3592],seed[2892],seed[2549],seed[357],seed[3595],seed[2116],seed[3849],seed[4078],seed[3354],seed[3399],seed[3079],seed[3395],seed[1934],seed[1170],seed[476],seed[3167],seed[2014],seed[2335],seed[3631],seed[600],seed[2540],seed[762],seed[3701],seed[2628],seed[1080],seed[478],seed[3922],seed[995],seed[1491],seed[3281],seed[553],seed[403],seed[127],seed[2275],seed[142],seed[364],seed[557],seed[3656],seed[2931],seed[3301],seed[3424],seed[3345],seed[2257],seed[773],seed[4012],seed[2174],seed[3068],seed[669],seed[1580],seed[3459],seed[163],seed[2409],seed[2278],seed[1777],seed[175],seed[2020],seed[3276],seed[2205],seed[3714],seed[3332],seed[3670],seed[1890],seed[2692],seed[1802],seed[463],seed[1877],seed[1878],seed[1701],seed[1859],seed[3435],seed[800],seed[1751],seed[3507],seed[3778],seed[4054],seed[2770],seed[1678],seed[1953],seed[1088],seed[224],seed[1728],seed[93],seed[3510],seed[970],seed[943],seed[1960],seed[3861],seed[2144],seed[3791],seed[2698],seed[798],seed[1224],seed[1514],seed[2066],seed[1686],seed[552],seed[3724],seed[3134],seed[867],seed[3420],seed[3935],seed[989],seed[3837],seed[64],seed[3007],seed[1],seed[529],seed[3425],seed[1882],seed[1196],seed[1898],seed[1068],seed[33],seed[4001],seed[2744],seed[2972],seed[444],seed[3540],seed[1444],seed[604],seed[1237],seed[1399],seed[2697],seed[2459],seed[1024],seed[3070],seed[1453],seed[3036],seed[3799],seed[173],seed[3763],seed[1557],seed[1419],seed[1570],seed[427],seed[1576],seed[2858],seed[1346],seed[2049],seed[3173],seed[2957],seed[473],seed[3503],seed[1706],seed[1526],seed[2869],seed[1033],seed[3066],seed[1427],seed[2838],seed[2168],seed[3076],seed[3965],seed[1300],seed[141],seed[741],seed[481],seed[2211],seed[2681],seed[3862],seed[1879],seed[3216],seed[2620],seed[1530],seed[2835],seed[514],seed[3893],seed[1733],seed[1061],seed[523],seed[2287],seed[1273],seed[2141],seed[872],seed[1804],seed[707],seed[3741],seed[2576],seed[2075],seed[1001],seed[2255],seed[2994],seed[2176],seed[382],seed[2088],seed[1100],seed[828],seed[233],seed[4092],seed[1329],seed[176],seed[550],seed[1041],seed[810],seed[4068],seed[2898],seed[3423],seed[2526],seed[2962],seed[1162],seed[1966],seed[3973],seed[383],seed[1588],seed[2366],seed[3689],seed[261],seed[785],seed[3859],seed[3147],seed[1552],seed[3571],seed[595],seed[1026],seed[238],seed[3321],seed[3866],seed[3924],seed[2961],seed[2565],seed[3820],seed[1605],seed[2927],seed[2945],seed[3063],seed[3635],seed[721],seed[3773],seed[964],seed[665],seed[236],seed[3754],seed[2139],seed[499],seed[2473],seed[2851],seed[2552],seed[968],seed[2837],seed[1830],seed[2442],seed[1522],seed[132],seed[1214],seed[3191],seed[1967],seed[1164],seed[2774],seed[2352],seed[1973],seed[1173],seed[2153],seed[503],seed[939],seed[3311],seed[2845],seed[2371],seed[3515],seed[3855],seed[2397],seed[1417],seed[3275],seed[3499],seed[4048],seed[578],seed[1543],seed[740],seed[873],seed[1999],seed[2166],seed[2805],seed[1025],seed[323],seed[3337],seed[3702],seed[645],seed[2467],seed[2407],seed[2820],seed[577],seed[1542],seed[3810],seed[2990],seed[461],seed[1321],seed[1398],seed[1904],seed[2312],seed[2334],seed[3552],seed[2114],seed[3449],seed[516],seed[2329],seed[2660],seed[3168],seed[256],seed[1203],seed[2795],seed[506],seed[276],seed[3159],seed[2133],seed[3180],seed[1320],seed[2694],seed[1141],seed[2358],seed[2923],seed[3790],seed[1547],seed[2776],seed[3721],seed[3673],seed[3272],seed[370],seed[3610],seed[1148],seed[2615],seed[2699],seed[2758],seed[3726],seed[3158],seed[753],seed[1910],seed[3383],seed[1867],seed[2500],seed[2484],seed[1902],seed[2353],seed[4084],seed[1157],seed[539],seed[3394],seed[3649],seed[3666],seed[3389],seed[3985],seed[733],seed[1045],seed[21],seed[2582],seed[2223],seed[3522],seed[1714],seed[3366],seed[1225],seed[106],seed[935],seed[1748],seed[1537],seed[2354],seed[1793],seed[1248],seed[3011],seed[381],seed[1950],seed[861],seed[3217],seed[1883],seed[691],seed[839],seed[1190],seed[3848],seed[1689],seed[1191],seed[2388],seed[1690],seed[3693],seed[3479],seed[484],seed[3440],seed[3439],seed[3351],seed[1497],seed[2965],seed[559],seed[1510],seed[2992],seed[2336],seed[3986],seed[1702],seed[1382],seed[1886],seed[1469],seed[3218],seed[1452],seed[2557],seed[1870],seed[833],seed[1594],seed[482],seed[1445],seed[2344],seed[2310],seed[2045],seed[2512],seed[1307],seed[771],seed[3995],seed[1246],seed[2064],seed[3981],seed[796],seed[3713],seed[2571],seed[2621],seed[1769],seed[2590],seed[3876],seed[541],seed[868],seed[1070],seed[2149],seed[2847],seed[643],seed[4034],seed[2855],seed[1663],seed[3761],seed[3264],seed[318],seed[254],seed[213],seed[3358],seed[2476],seed[3725],seed[3787],seed[3511],seed[1211],seed[290],seed[3190],seed[489],seed[3756],seed[1880],seed[3145],seed[1659],seed[3512],seed[2806],seed[623],seed[592],seed[3172],seed[1117],seed[3581],seed[3436],seed[6],seed[1128],seed[2000],seed[3867],seed[2475],seed[2417],seed[3452],seed[2213],seed[2238],seed[1351],seed[3177],seed[915],seed[3333],seed[793],seed[587],seed[1603],seed[328],seed[2986],seed[1433],seed[1139],seed[1528],seed[2362],seed[957],seed[1501],seed[634],seed[3080],seed[1597],seed[2902],seed[1838],seed[2784],seed[20],seed[1865],seed[954],seed[548],seed[3716],seed[2303],seed[2588],seed[2634],seed[3115],seed[4013],seed[299],seed[2914],seed[4027],seed[1242],seed[2625],seed[3968],seed[2186],seed[2741],seed[479],seed[765],seed[1740],seed[1638],seed[2458],seed[1513],seed[1106],seed[648],seed[752],seed[3304],seed[3643],seed[2731],seed[2293],seed[1764],seed[1948],seed[2513],seed[2239],seed[2330],seed[3987],seed[3470],seed[1945],seed[3938],seed[2299],seed[2530],seed[1483],seed[1016],seed[2963],seed[2259],seed[1695],seed[4085],seed[1310],seed[2005],seed[3586],seed[1301],seed[2393],seed[893],seed[3071],seed[3789],seed[1863],seed[3890],seed[678],seed[744],seed[186],seed[319],seed[2323],seed[248],seed[2740],seed[120],seed[2403],seed[1642],seed[1636],seed[2155],seed[53],seed[73],seed[4041],seed[2097],seed[321],seed[540],seed[3003],seed[2651],seed[2844],seed[629],seed[2118],seed[2261],seed[809],seed[681],seed[1050],seed[895],seed[2607],seed[180],seed[2522],seed[29],seed[2750],seed[1335],seed[714],seed[3877],seed[2534],seed[63],seed[985],seed[818],seed[422],seed[3398],seed[2089],seed[2870],seed[2055],seed[1165],seed[3472],seed[3513],seed[1700],seed[1442],seed[3871],seed[3710],seed[1736],seed[842],seed[1896],seed[1352],seed[3530],seed[3232],seed[2111],seed[360],seed[3161],seed[823],seed[3630],seed[3490],seed[2194],seed[27],seed[509],seed[2180],seed[857],seed[367],seed[1574],seed[2214],seed[4058],seed[3842],seed[615],seed[1517],seed[3469],seed[3139],seed[1463],seed[2886],seed[2337],seed[1258],seed[3315],seed[136],seed[153],seed[2626],seed[1030],seed[1272],seed[2480],seed[313],seed[2463],seed[204],seed[565],seed[2829],seed[2742],seed[1076],seed[3591],seed[3361],seed[1874],seed[3160],seed[2283],seed[3647],seed[3455],seed[3213],seed[2306],seed[2678],seed[3092],seed[2777],seed[631],seed[96],seed[3342],seed[2162],seed[1441],seed[1012],seed[86],seed[2722],seed[341],seed[1791],seed[4003],seed[2215],seed[3750],seed[981],seed[162],seed[1087],seed[2209],seed[3900],seed[925],seed[55],seed[3528],seed[764],seed[3138],seed[649],seed[2202],seed[3331],seed[3223],seed[2233],seed[3025],seed[1350],seed[212],seed[2224],seed[2217],seed[3075],seed[2779],seed[2908],seed[258],seed[3257],seed[2394],seed[1311],seed[1726],seed[3294],seed[3340],seed[1872],seed[3114],seed[1641],seed[3121],seed[1306],seed[2716],seed[3846],seed[220],seed[2591],seed[269],seed[1954],seed[2496],seed[1653],seed[1357],seed[1048],seed[152],seed[3157],seed[1851],seed[2443],seed[3578],seed[1620],seed[2433],seed[1541],seed[808],seed[2826],seed[1651],seed[457],seed[3429],seed[2083],seed[2989],seed[2984],seed[1795],seed[234],seed[1402],seed[3650],seed[1199],seed[2754],seed[1850],seed[1334],seed[1718],seed[4024],seed[3185],seed[3879],seed[889],seed[1102],seed[50],seed[1515],seed[1734],seed[502],seed[3916],seed[651],seed[449],seed[3770],seed[974],seed[2262],seed[464],seed[1852],seed[982],seed[293],seed[3776],seed[513],seed[3950],seed[339],seed[26],seed[3764],seed[3244],seed[2786],seed[1573],seed[3736],seed[2932],seed[1676],seed[3963],seed[2482],seed[5],seed[3461],seed[1280],seed[1057],seed[3894],seed[2551],seed[736],seed[245],seed[3197],seed[2712],seed[3887],seed[1941],seed[920],seed[2926],seed[2996],seed[2884],seed[3280],seed[480],seed[528],seed[1712],seed[2737],seed[1683],seed[992],seed[698],seed[1397],seed[3732],seed[705],seed[3427],seed[1741],seed[354],seed[2241],seed[1575],seed[2680],seed[78],seed[2947],seed[3830],seed[2816],seed[2419],seed[1823],seed[3579],seed[2343],seed[3585],seed[2675],seed[3590],seed[515],seed[3187],seed[3060],seed[4009],seed[3942],seed[3840],seed[3806],seed[47],seed[30],seed[668],seed[3538],seed[3816],seed[716],seed[4086],seed[2135],seed[1285],seed[2514],seed[609],seed[2956],seed[3006],seed[1027],seed[184],seed[2519],seed[1363],seed[690],seed[419],seed[410],seed[2631],seed[599],seed[1449],seed[1053],seed[1021],seed[2210],seed[2661],seed[1884],seed[1275],seed[3671],seed[961],seed[100],seed[551],seed[3672],seed[4069],seed[3795],seed[104],seed[2528],seed[2646],seed[3230],seed[1822],seed[2120],seed[447],seed[2663],seed[468],seed[3417],seed[3203],seed[2974],seed[803],seed[438],seed[61],seed[3874],seed[3542],seed[2558],seed[1145],seed[1496],seed[955],seed[3444],seed[3569],seed[537],seed[462],seed[1460],seed[1118],seed[4056],seed[2719],seed[43],seed[2325],seed[2225],seed[619],seed[1215],seed[168],seed[3829],seed[2943],seed[2359],seed[3660],seed[1832],seed[3782],seed[3823],seed[3574],seed[1719],seed[415],seed[2367],seed[445],seed[704],seed[3181],seed[1015],seed[3206],seed[3289],seed[1368],seed[260],seed[3651],seed[3988],seed[34],seed[2346],seed[945],seed[190],seed[3905],seed[672],seed[3371],seed[3551],seed[3105],seed[997],seed[2815],seed[126],seed[3629],seed[998],seed[1425],seed[198],seed[2372],seed[2728],seed[3314],seed[3313],seed[1790],seed[3027],seed[973],seed[3090],seed[567],seed[2599],seed[797],seed[1189],seed[4077],seed[237],seed[726],seed[2052],seed[2733],seed[784],seed[1161],seed[1342],seed[3722],seed[1333],seed[241],seed[642],seed[1339],seed[2331],seed[2587],seed[2054],seed[1341],seed[1479],seed[1564],seed[1824],seed[2955],seed[3558],seed[2801],seed[2044],seed[3653],seed[202],seed[286],seed[3271],seed[3221],seed[3214],seed[1049],seed[790],seed[310],seed[1366],seed[3299],seed[2445],seed[3664],seed[1648],seed[3184],seed[2515],seed[1315],seed[2253],seed[349],seed[196],seed[231],seed[2987],seed[3792],seed[3409],seed[1018],seed[2497],seed[3700],seed[3723],seed[2667],seed[3970],seed[3914],seed[3169],seed[1410],seed[44],seed[2307],seed[927],seed[646],seed[558],seed[70],seed[1956],seed[3194],seed[336],seed[340],seed[368],seed[1707],seed[4065],seed[2189],seed[3777],seed[1055],seed[2086],seed[3245],seed[743],seed[2148],seed[3428],seed[792],seed[4011],seed[284],seed[3051],seed[1722],seed[2041],seed[1287],seed[944],seed[1362],seed[262],seed[2669],seed[1652],seed[3753],seed[1328],seed[2494],seed[622],seed[1168],seed[3086],seed[779],seed[2804],seed[2852],seed[1197],seed[879],seed[2933],seed[2903],seed[110],seed[1847],seed[782],seed[1876],seed[3305],seed[1598],seed[1418],seed[1426],seed[2332],seed[3231],seed[2108],seed[3917],seed[4031],seed[1658],seed[1939],seed[3962],seed[477],seed[11],seed[2853],seed[1127],seed[2471],seed[434],seed[1174],seed[852],seed[1308],seed[388],seed[1798],seed[582],seed[712],seed[49],seed[696],seed[3235],seed[1082],seed[3433],seed[3162],seed[1861],seed[366],seed[3881],seed[2944],seed[2517],seed[501],seed[3620],seed[244],seed[3128],seed[2110],seed[1871],seed[2489],seed[3555],seed[2079],seed[3593],seed[1279],seed[3596],seed[3493],seed[3042],seed[3797],seed[2474],seed[1042],seed[1679],seed[1421],seed[888],seed[2887],seed[2199],seed[3899],seed[4029],seed[3239],seed[1922],seed[3918],seed[2501],seed[1912],seed[475],seed[887],seed[3587],seed[208],seed[1464],seed[2095],seed[2717],seed[1908],seed[2734],seed[2232],seed[2434],seed[2015],seed[2381],seed[1775],seed[433],seed[1729],seed[2308],seed[3734],seed[3925],seed[3317],seed[4021],seed[947],seed[374],seed[1354],seed[3378],seed[2430],seed[2314],seed[606],seed[183],seed[1038],seed[1099],seed[80],seed[1782],seed[3329],seed[996],seed[2830],seed[2521],seed[2400],seed[3293],seed[2601],seed[870],seed[1457],seed[3041],seed[3527],seed[2511],seed[2068],seed[2121],seed[2564],seed[1807],seed[3016],seed[802],seed[3083],seed[1458],seed[279],seed[2899],seed[693],seed[2305],seed[452],seed[848],seed[3376],seed[3597],seed[3544],seed[824],seed[1104],seed[218],seed[1812],seed[1438],seed[2585],seed[16],seed[1487],seed[2876],seed[1195],seed[1800],seed[1212],seed[1202],seed[265],seed[1098],seed[3944],seed[255],seed[684],seed[1493],seed[3055],seed[3397],seed[2297],seed[1788],seed[4051],seed[266],seed[1240],seed[1688],seed[1944],seed[3854],seed[440],seed[2860],seed[342],seed[2438],seed[2469],seed[376],seed[2012],seed[1052],seed[1713],seed[134],seed[1256],seed[906],seed[2439],seed[414],seed[1836],seed[904],seed[3719],seed[3010],seed[2539],seed[1602],seed[2589],seed[3316],seed[1993],seed[2460],seed[160],seed[2405],seed[3807],seed[3343],seed[3065],seed[564],seed[1596],seed[250],seed[103],seed[2242],seed[1423],seed[4023],seed[2190],seed[264],seed[3116],seed[1336],seed[1490],seed[486],seed[2247],seed[453],seed[2156],seed[825],seed[2817],seed[1579],seed[1090],seed[2819],seed[2119],seed[3688],seed[846],seed[3793],seed[3869],seed[3155],seed[4040],seed[3652],seed[3897],seed[283],seed[3910],seed[2873],seed[3783],seed[3765],seed[821],seed[1465],seed[2723],seed[3103],seed[3589],seed[962],seed[2037],seed[2413],seed[1732],seed[2708],seed[1855],seed[3766],seed[2132],seed[3934],seed[15],seed[1373],seed[2435],seed[3390],seed[3568],seed[1276],seed[3338],seed[1585],seed[533],seed[3641],seed[1554],seed[1407],seed[320],seed[470],seed[835],seed[1619],seed[1892],seed[3393],seed[3309],seed[3062],seed[2848],seed[3432],seed[3038],seed[3094],seed[2270],seed[1796],seed[3437],seed[3211],seed[2755],seed[4087],seed[1370],seed[1304],seed[676],seed[1601],seed[3932],seed[851],seed[3457],seed[1503],seed[3384],seed[3325],seed[3863],seed[3467],seed[48],seed[1123],seed[94],seed[1432],seed[267],seed[54],seed[1002],seed[2709],seed[1192],seed[3911],seed[2129],seed[884],seed[1685],seed[2854],seed[795],seed[4049],seed[2940],seed[2],seed[2046],seed[739],seed[2462],seed[929],seed[3248],seed[1909],seed[206],seed[3500],seed[1365],seed[2245],seed[2374],seed[2103],seed[1481],seed[330],seed[2277],seed[2207],seed[1935],seed[1744],seed[3502],seed[4075],seed[2533],seed[3901],seed[3561],seed[3892],seed[2465],seed[2715],seed[2100],seed[1825],seed[695],seed[841],seed[3994],seed[3273],seed[2237],seed[2548],seed[826],seed[426],seed[3506],seed[1520],seed[1209],seed[692],seed[1622],seed[1784],seed[3403],seed[2197],seed[2968],seed[277],seed[1887],seed[2798],seed[727],seed[1089],seed[2952],seed[3445],seed[3712],seed[2195],seed[1618],seed[2527],seed[2605],seed[3012],seed[88],seed[498],seed[3550],seed[2743],seed[614],seed[1862],seed[3687],seed[385],seed[2971],seed[2383],seed[1376],seed[3339],seed[677],seed[2043],seed[2432],seed[898],seed[657],seed[2633],seed[2609],seed[1931],seed[3612],seed[3501],seed[2013],seed[1292],seed[2017],seed[2090],seed[287],seed[3902],seed[3170],seed[1096],seed[2415],seed[1241],seed[3410],seed[1151],seed[1660],seed[3441],seed[610],seed[1593],seed[273],seed[778],seed[1155],seed[4037],seed[2939],seed[3553],seed[538],seed[2333],seed[750],seed[3246],seed[2595],seed[131],seed[2597],seed[101],seed[2254],seed[1271],seed[3456],seed[1232],seed[554],seed[2904],seed[3415],seed[1894],seed[2928],seed[862],seed[1779],seed[2641],seed[2790],seed[3563],seed[4063],seed[2524],seed[775],seed[2724],seed[1581],seed[118],seed[3302],seed[1578],seed[1738],seed[2127],seed[2175],seed[956],seed[612],seed[1044],seed[226],seed[2686],seed[1889],seed[1929],seed[1994],seed[2897],seed[2488],seed[3801],seed[1727],seed[2654],seed[459],seed[2577],seed[2117],seed[1152],seed[1138],seed[191],seed[1617],seed[1439],seed[3802],seed[3600],seed[111],seed[517],seed[10],seed[1381],seed[1325],seed[1182],seed[3192],seed[2092],seed[3885],seed[1008],seed[2137],seed[880],seed[3295],seed[923],seed[2655],seed[701],seed[1509],seed[863],seed[1097],seed[1817],seed[2154],seed[3448],seed[1236],seed[3781],seed[3744],seed[2556],seed[4081],seed[257],seed[2840],seed[2814],seed[3023],seed[3800],seed[1286],seed[1175],seed[4033],seed[546],seed[4039],seed[2248],seed[3960],seed[3233],seed[3533],seed[2802],seed[3150],seed[979],seed[1468],seed[670],seed[734],seed[154],seed[983],seed[1422],seed[3207],seed[1109],seed[1819],seed[1019],seed[1416],seed[1746],seed[3269],seed[2762],seed[1259],seed[2685],seed[1229],seed[1942],seed[441],seed[3225],seed[2993],seed[2377],seed[2690],seed[1014],seed[439],seed[2282],seed[2035],seed[192],seed[1348],seed[3357],seed[535],seed[3268],seed[799],seed[2326],seed[1961],seed[1217],seed[259],seed[2711],seed[3200],seed[3179],seed[2418],seed[2219],seed[4072],seed[3431],seed[2146],seed[2818],seed[4032],seed[3780],seed[292],seed[1697],seed[1078],seed[2510],seed[334],seed[22],seed[1749],seed[738],seed[1661],seed[2954],seed[3692],seed[3904],seed[3263],seed[518],seed[4036],seed[3992],seed[2427],seed[1955],seed[3262],seed[2266],seed[2437],seed[2547],seed[2905],seed[2662],seed[129],seed[3048],seed[3064],seed[413],seed[2423],seed[2689],seed[1213],seed[3040],seed[4042],seed[2112],seed[4005],seed[3704],seed[2696],seed[1525],seed[2682],seed[3084],seed[3858],seed[1972],seed[1171],seed[4076],seed[2378],seed[1101],seed[2385],seed[2760],seed[3737],seed[1343],seed[0],seed[3237],seed[1226],seed[2436],seed[2264],seed[1924],seed[2793],seed[2159],seed[2614],seed[2102],seed[2051],seed[3541],seed[1251],seed[92],seed[17],seed[952],seed[1112],seed[1533],seed[327],seed[3727],seed[758],seed[2039],seed[1773],seed[2229],seed[3525],seed[3146],seed[1958],seed[3001],seed[975],seed[3570],seed[4070],seed[246],seed[1551],seed[859],seed[210],seed[3755],seed[2322],seed[1461],seed[3696],seed[4061],seed[1230],seed[1845],seed[1456],seed[536],seed[371],seed[2392],seed[1377],seed[3481],seed[530],seed[195],seed[280],seed[2763],seed[656],seed[2752],seed[1281],seed[2613],seed[4094],seed[1628],seed[1521],seed[156],seed[338],seed[3270],seed[2543],seed[1081],seed[1755],seed[3201],seed[3183],seed[2263],seed[2866],seed[3821],seed[2291],seed[2649],seed[1115],seed[2398],seed[2574],seed[855],seed[2502],seed[768],seed[1981],seed[124],seed[2252],seed[2532],seed[1066],seed[1404],seed[1201],seed[329],seed[1186],seed[2505],seed[2778],seed[3627],seed[2583],seed[2768],seed[1974],seed[487],seed[630],seed[2748],seed[2594],seed[408],seed[140],seed[1634],seed[3749],seed[1114],seed[1359],seed[324],seed[159],seed[3101],seed[659],seed[2258],seed[1331],seed[2856],seed[3222],seed[1849],seed[3303],seed[1947],seed[1621],seed[2338],seed[85],seed[840],seed[932],seed[1868],seed[2650],seed[358],seed[827],seed[1144],seed[1977],seed[3891],seed[3564],seed[625],seed[4059],seed[2629],seed[1111],seed[2324],seed[1895],seed[2379],seed[3974],seed[1508],seed[229],seed[628],seed[38],seed[3531],seed[2756],seed[1703],seed[387],seed[1126],seed[1899],seed[3081],seed[2289],seed[2216],seed[8],seed[1997],seed[3067],seed[2773],seed[3004],seed[3348],seed[421],seed[1682],seed[3405],seed[3928],seed[405],seed[757],seed[3662],seed[189],seed[723],seed[3059],seed[65],seed[1649],seed[2455],seed[1250],seed[1347],seed[1265],seed[2976],seed[3768],seed[2163],seed[3053],seed[3199],seed[667],seed[3095],seed[418],seed[1293],seed[337],seed[1472],seed[2880],seed[3638],seed[1208],seed[2274],seed[519],seed[3381],seed[3069],seed[3226],seed[3484],seed[2783],seed[885],seed[1235],seed[972],seed[3024],seed[1047],seed[3240],seed[2647],seed[1615],seed[3955],seed[46],seed[2537],seed[251],seed[2152],seed[451],seed[1831],seed[3093],seed[918],seed[2827]}),
        .cross_prob(cross_prob),
        .codeword(codeword4),
        .received(received4)
        );
    
    bsc bsc5(
        .clk(clk),
        .reset(reset),
        .seed({seed[2337],seed[1934],seed[1406],seed[2097],seed[1209],seed[623],seed[2156],seed[2843],seed[3321],seed[2529],seed[1042],seed[617],seed[227],seed[636],seed[2499],seed[2679],seed[396],seed[882],seed[2662],seed[3776],seed[3946],seed[3628],seed[1082],seed[3061],seed[1675],seed[3639],seed[2907],seed[990],seed[2563],seed[3837],seed[1030],seed[3616],seed[3144],seed[1670],seed[2038],seed[2865],seed[2167],seed[3093],seed[3733],seed[3081],seed[1625],seed[3676],seed[3025],seed[3454],seed[484],seed[3100],seed[2113],seed[1129],seed[715],seed[3045],seed[1328],seed[1038],seed[2225],seed[2164],seed[3929],seed[3147],seed[1172],seed[945],seed[3720],seed[1390],seed[278],seed[3356],seed[3878],seed[651],seed[3413],seed[933],seed[1352],seed[3752],seed[3692],seed[2240],seed[2789],seed[112],seed[1431],seed[3654],seed[2596],seed[621],seed[2311],seed[3652],seed[2218],seed[2883],seed[3274],seed[1252],seed[2964],seed[2166],seed[1800],seed[372],seed[2356],seed[521],seed[3175],seed[3912],seed[4022],seed[1037],seed[2944],seed[3255],seed[2953],seed[1467],seed[2176],seed[2556],seed[1768],seed[1512],seed[3031],seed[123],seed[837],seed[3779],seed[1210],seed[902],seed[2895],seed[1391],seed[738],seed[2109],seed[1114],seed[821],seed[1147],seed[2458],seed[972],seed[1740],seed[3816],seed[3780],seed[2009],seed[3207],seed[813],seed[81],seed[644],seed[1191],seed[1382],seed[3458],seed[1417],seed[3542],seed[3861],seed[1557],seed[3462],seed[1614],seed[3990],seed[1872],seed[3782],seed[2005],seed[3334],seed[1330],seed[384],seed[3104],seed[4063],seed[734],seed[3787],seed[512],seed[3243],seed[2608],seed[1908],seed[2383],seed[1485],seed[236],seed[53],seed[1696],seed[576],seed[2373],seed[1663],seed[1763],seed[3727],seed[1664],seed[1769],seed[452],seed[113],seed[2721],seed[3027],seed[13],seed[3544],seed[3532],seed[3993],seed[1795],seed[3171],seed[3739],seed[3295],seed[2191],seed[539],seed[2532],seed[2574],seed[3710],seed[2346],seed[475],seed[2763],seed[489],seed[3869],seed[1111],seed[591],seed[2654],seed[72],seed[733],seed[300],seed[1651],seed[3392],seed[936],seed[2619],seed[987],seed[662],seed[2444],seed[3037],seed[1597],seed[3564],seed[2023],seed[3914],seed[1883],seed[420],seed[3693],seed[1238],seed[947],seed[3264],seed[2727],seed[4046],seed[2677],seed[3999],seed[811],seed[1929],seed[3862],seed[3822],seed[3437],seed[2012],seed[1548],seed[2811],seed[2650],seed[1452],seed[1949],seed[3279],seed[1353],seed[2448],seed[3358],seed[3699],seed[1764],seed[2273],seed[732],seed[2836],seed[2110],seed[30],seed[391],seed[1882],seed[3096],seed[1412],seed[3698],seed[3103],seed[1376],seed[2316],seed[216],seed[96],seed[2745],seed[142],seed[602],seed[2586],seed[2561],seed[1277],seed[307],seed[3870],seed[3026],seed[3823],seed[2548],seed[2293],seed[2613],seed[1263],seed[2967],seed[3339],seed[741],seed[1011],seed[3820],seed[3346],seed[2050],seed[543],seed[2656],seed[1954],seed[1781],seed[3051],seed[41],seed[2],seed[831],seed[11],seed[3700],seed[3677],seed[1013],seed[1043],seed[2090],seed[509],seed[347],seed[2894],seed[2011],seed[2231],seed[2801],seed[3411],seed[1688],seed[1427],seed[867],seed[298],seed[3706],seed[725],seed[329],seed[1257],seed[1531],seed[373],seed[3017],seed[1225],seed[1092],seed[1824],seed[706],seed[542],seed[2436],seed[27],seed[736],seed[879],seed[392],seed[2220],seed[1308],seed[2179],seed[1091],seed[2234],seed[1870],seed[3962],seed[2454],seed[1451],seed[2208],seed[1957],seed[3432],seed[3245],seed[1060],seed[3858],seed[1588],seed[2777],seed[1628],seed[1029],seed[3211],seed[1283],seed[150],seed[1141],seed[4059],seed[3079],seed[116],seed[845],seed[1259],seed[3040],seed[4029],seed[1154],seed[3403],seed[3593],seed[2972],seed[1297],seed[352],seed[2196],seed[1912],seed[2425],seed[2765],seed[3755],seed[1359],seed[1018],seed[359],seed[2204],seed[1735],seed[3927],seed[153],seed[787],seed[4048],seed[3748],seed[2517],seed[3164],seed[4068],seed[33],seed[3716],seed[4004],seed[2950],seed[795],seed[2708],seed[1344],seed[1443],seed[2267],seed[1317],seed[1070],seed[3267],seed[1533],seed[4028],seed[2615],seed[2370],seed[1095],seed[2392],seed[2036],seed[3817],seed[1522],seed[1930],seed[3498],seed[3934],seed[754],seed[2987],seed[2739],seed[642],seed[1838],seed[331],seed[2916],seed[1404],seed[518],seed[1933],seed[3029],seed[1349],seed[3401],seed[628],seed[680],seed[763],seed[1447],seed[3224],seed[1160],seed[2887],seed[2636],seed[3886],seed[1939],seed[469],seed[1545],seed[3890],seed[3673],seed[1825],seed[4067],seed[2978],seed[1757],seed[1266],seed[2527],seed[344],seed[2158],seed[136],seed[917],seed[78],seed[403],seed[2178],seed[408],seed[2882],seed[10],seed[2354],seed[2086],seed[3873],seed[69],seed[529],seed[701],seed[208],seed[3501],seed[34],seed[2531],seed[2287],seed[3249],seed[1026],seed[3888],seed[789],seed[792],seed[2157],seed[4018],seed[2378],seed[1798],seed[633],seed[2457],seed[2500],seed[3278],seed[435],seed[793],seed[1459],seed[526],seed[2989],seed[525],seed[209],seed[3588],seed[3907],seed[851],seed[429],seed[1902],seed[3519],seed[1102],seed[1839],seed[908],seed[2889],seed[1604],seed[1186],seed[3032],seed[2886],seed[2075],seed[3333],seed[107],seed[188],seed[1881],seed[1595],seed[324],seed[3713],seed[1040],seed[618],seed[886],seed[575],seed[211],seed[131],seed[2081],seed[3416],seed[3536],seed[67],seed[993],seed[961],seed[3611],seed[3814],seed[2830],seed[530],seed[196],seed[3766],seed[1988],seed[2728],seed[2984],seed[3859],seed[1059],seed[3439],seed[3304],seed[531],seed[1906],seed[2798],seed[1674],seed[2908],seed[3145],seed[678],seed[2911],seed[1634],seed[3273],seed[1851],seed[681],seed[1446],seed[3417],seed[2736],seed[3374],seed[2439],seed[3500],seed[1239],seed[466],seed[1201],seed[742],seed[1471],seed[2228],seed[629],seed[1190],seed[3894],seed[1931],seed[957],seed[2121],seed[1559],seed[645],seed[3446],seed[1363],seed[3453],seed[1943],seed[2324],seed[968],seed[1233],seed[1613],seed[3470],seed[2520],seed[3138],seed[3496],seed[1525],seed[3599],seed[747],seed[1206],seed[288],seed[256],seed[3441],seed[1509],seed[140],seed[1249],seed[2014],seed[2847],seed[2623],seed[1304],seed[520],seed[3572],seed[3734],seed[1842],seed[2330],seed[2526],seed[1341],seed[1272],seed[3187],seed[2415],seed[2738],seed[230],seed[1395],seed[1987],seed[3041],seed[467],seed[684],seed[105],seed[12],seed[3158],seed[303],seed[1913],seed[294],seed[3595],seed[3580],seed[3],seed[951],seed[3574],seed[2575],seed[1243],seed[1486],seed[1834],seed[3003],seed[2275],seed[2091],seed[816],seed[14],seed[339],seed[1847],seed[2203],seed[1647],seed[2676],seed[3113],seed[523],seed[1397],seed[3798],seed[2729],seed[2602],seed[2923],seed[3913],seed[1985],seed[1563],seed[2408],seed[4001],seed[1492],seed[941],seed[1106],seed[190],seed[4033],seed[1130],seed[1547],seed[551],seed[277],seed[1889],seed[2338],seed[2667],seed[900],seed[1997],seed[219],seed[312],seed[1136],seed[3456],seed[1739],seed[2928],seed[427],seed[1966],seed[2332],seed[267],seed[603],seed[2379],seed[167],seed[594],seed[1150],seed[3343],seed[519],seed[1683],seed[1978],seed[2760],seed[2162],seed[2404],seed[2762],seed[2835],seed[1333],seed[280],seed[2029],seed[3575],seed[1510],seed[953],seed[4088],seed[2302],seed[438],seed[4065],seed[2771],seed[1950],seed[343],seed[2349],seed[3603],seed[712],seed[3989],seed[1762],seed[1032],seed[18],seed[977],seed[1483],seed[3420],seed[3924],seed[315],seed[3825],seed[2595],seed[1846],seed[2910],seed[301],seed[1741],seed[2512],seed[2455],seed[859],seed[1806],seed[3657],seed[1539],seed[895],seed[2295],seed[2319],seed[2783],seed[1594],seed[3265],seed[1320],seed[3773],seed[3302],seed[3597],seed[3645],seed[1526],seed[2694],seed[2185],seed[1074],seed[4011],seed[1843],seed[2306],seed[989],seed[2871],seed[2627],seed[1809],seed[3505],seed[2549],seed[685],seed[599],seed[2990],seed[973],seed[2852],seed[95],seed[3561],seed[2460],seed[3976],seed[173],seed[36],seed[1515],seed[1265],seed[370],seed[2732],seed[2219],seed[812],seed[2447],seed[597],seed[2312],seed[260],seed[2441],seed[1161],seed[1462],seed[2993],seed[627],seed[3303],seed[814],seed[1294],seed[1875],seed[3843],seed[1714],seed[1772],seed[3436],seed[434],seed[1529],seed[3445],seed[4003],seed[2135],seed[3694],seed[1876],seed[2484],seed[2027],seed[2296],seed[1151],seed[2700],seed[753],seed[16],seed[3757],seed[2860],seed[1873],seed[2599],seed[1008],seed[1401],seed[3162],seed[1558],seed[2045],seed[1168],seed[2122],seed[975],seed[3393],seed[829],seed[1569],seed[2340],seed[3877],seed[616],seed[3384],seed[515],seed[2276],seed[3076],seed[1478],seed[4053],seed[1561],seed[1436],seed[2400],seed[3370],seed[1377],seed[2658],seed[2125],seed[1700],seed[2797],seed[3534],seed[317],seed[1699],seed[3607],seed[1895],seed[3939],seed[1188],seed[2977],seed[1226],seed[892],seed[3805],seed[316],seed[841],seed[871],seed[120],seed[2107],seed[3804],seed[2968],seed[746],seed[1274],seed[562],seed[117],seed[2854],seed[1348],seed[1612],seed[266],seed[868],seed[3360],seed[1835],seed[2969],seed[415],seed[2335],seed[547],seed[2689],seed[929],seed[3231],seed[1915],seed[3975],seed[2069],seed[1468],seed[456],seed[1830],seed[2813],seed[3533],seed[1463],seed[3233],seed[25],seed[1223],seed[440],seed[728],seed[411],seed[3788],seed[3553],seed[1244],seed[1474],seed[3083],seed[3627],seed[2453],seed[3925],seed[3021],seed[2022],seed[943],seed[985],seed[2190],seed[2872],seed[1788],seed[2795],seed[561],seed[827],seed[2681],seed[3022],seed[3062],seed[463],seed[3560],seed[1543],seed[302],seed[1110],seed[2628],seed[253],seed[1606],seed[1598],seed[1291],seed[788],seed[3653],seed[103],seed[4056],seed[3316],seed[3524],seed[3214],seed[2937],seed[2384],seed[306],seed[2181],seed[2412],seed[528],seed[3452],seed[43],seed[3831],seed[1019],seed[3151],seed[2539],seed[3306],seed[1442],seed[2072],seed[308],seed[2361],seed[44],seed[1626],seed[1068],seed[3232],seed[2980],seed[2294],seed[1221],seed[1975],seed[3320],seed[1012],seed[815],seed[3090],seed[1910],seed[2470],seed[579],seed[1343],seed[3209],seed[919],seed[1437],seed[3291],seed[1425],seed[174],seed[1952],seed[2868],seed[830],seed[2901],seed[3661],seed[590],seed[3218],seed[222],seed[3863],seed[2469],seed[2272],seed[735],seed[220],seed[2202],seed[3849],seed[3717],seed[2226],seed[1925],seed[3997],seed[1083],seed[1645],seed[675],seed[283],seed[844],seed[1681],seed[1819],seed[1938],seed[3827],seed[2982],seed[2318],seed[202],seed[3153],seed[2194],seed[2345],seed[273],seed[4015],seed[3821],seed[3747],seed[1560],seed[2610],seed[3590],seed[2925],seed[35],seed[3967],seed[1833],seed[233],seed[3811],seed[2479],seed[265],seed[803],seed[412],seed[3577],seed[1702],seed[1665],seed[2503],seed[444],seed[3922],seed[544],seed[2921],seed[905],seed[2633],seed[1776],seed[3485],seed[1310],seed[2971],seed[883],seed[1789],seed[4002],seed[2711],seed[2853],seed[175],seed[394],seed[1067],seed[2747],seed[1815],seed[1386],seed[3053],seed[3951],seed[171],seed[3292],seed[3495],seed[2101],seed[2104],seed[2954],seed[1078],seed[2433],seed[2616],seed[2806],seed[1305],seed[3228],seed[2651],seed[2594],seed[2822],seed[834],seed[620],seed[1995],seed[58],seed[2951],seed[1046],seed[1637],seed[1254],seed[1980],seed[3484],seed[1045],seed[1517],seed[39],seed[1077],seed[2848],seed[3276],seed[2037],seed[3486],seed[3672],seed[791],seed[2334],seed[181],seed[571],seed[3832],seed[1087],seed[1339],seed[1450],seed[3298],seed[3330],seed[3348],seed[1750],seed[2071],seed[3740],seed[1629],seed[672],seed[3902],seed[376],seed[1175],seed[3527],seed[655],seed[3957],seed[2932],seed[3014],seed[2170],seed[1361],seed[3425],seed[2111],seed[4066],seed[1063],seed[3647],seed[2067],seed[473],seed[4076],seed[799],seed[2857],seed[2252],seed[880],seed[1373],seed[3619],seed[3737],seed[2123],seed[3867],seed[3085],seed[221],seed[454],seed[2614],seed[102],seed[3404],seed[3891],seed[2592],seed[59],seed[566],seed[1421],seed[2945],seed[1648],seed[1234],seed[694],seed[3917],seed[1935],seed[1787],seed[2380],seed[3492],seed[4075],seed[311],seed[1718],seed[749],seed[45],seed[659],seed[2264],seed[3338],seed[2438],seed[138],seed[1156],seed[906],seed[1671],seed[3400],seed[2652],seed[2047],seed[364],seed[3082],seed[1192],seed[2829],seed[609],seed[619],seed[3736],seed[4077],seed[3389],seed[925],seed[1897],seed[1155],seed[3963],seed[739],seed[2746],seed[3034],seed[3613],seed[3691],seed[1752],seed[2348],seed[1023],seed[1942],seed[1917],seed[1860],seed[291],seed[2544],seed[564],seed[1241],seed[3714],seed[1643],seed[1736],seed[2501],seed[362],seed[3440],seed[205],seed[3379],seed[3764],seed[4034],seed[3852],seed[240],seed[3216],seed[3974],seed[3487],seed[3129],seed[481],seed[499],seed[3668],seed[3410],seed[305],seed[2618],seed[3357],seed[3217],seed[1774],seed[422],seed[1587],seed[1524],seed[313],seed[4085],seed[3636],seed[605],seed[1608],seed[1928],seed[1189],seed[2054],seed[3336],seed[3067],seed[1962],seed[1108],seed[1289],seed[3020],seed[3068],seed[2714],seed[1124],seed[2401],seed[3006],seed[3469],seed[3756],seed[2986],seed[4078],seed[1231],seed[2817],seed[1103],seed[1113],seed[607],seed[1396],seed[1368],seed[1242],seed[3666],seed[2118],seed[2748],seed[2959],seed[1213],seed[248],seed[3376],seed[3637],seed[3937],seed[3301],seed[4061],seed[166],seed[84],seed[3868],seed[1292],seed[3632],seed[3526],seed[580],seed[3172],seed[1378],seed[3133],seed[3194],seed[1552],seed[634],seed[955],seed[1687],seed[3464],seed[75],seed[2326],seed[121],seed[1281],seed[1355],seed[1017],seed[2686],seed[281],seed[3841],seed[836],seed[650],seed[2961],seed[1677],seed[3882],seed[1022],seed[2193],seed[2492],seed[432],seed[2612],seed[3378],seed[477],seed[2286],seed[3514],seed[1749],seed[660],seed[904],seed[3508],seed[3258],seed[2754],seed[2119],seed[262],seed[549],seed[3516],seed[1753],seed[3792],seed[3898],seed[3284],seed[326],seed[2182],seed[193],seed[360],seed[3846],seed[1465],seed[3406],seed[4019],seed[2692],seed[296],seed[2825],seed[1069],seed[805],seed[2581],seed[1163],seed[2973],seed[1907],seed[3328],seed[1250],seed[1432],seed[3537],seed[764],seed[1285],seed[1248],seed[3933],seed[2148],seed[2743],seed[237],seed[249],seed[1998],seed[1590],seed[1400],seed[3916],seed[2828],seed[1573],seed[2270],seed[1863],seed[3098],seed[1205],seed[3550],seed[2884],seed[322],seed[3540],seed[1521],seed[1593],seed[1801],seed[346],seed[48],seed[3159],seed[1454],seed[2976],seed[2502],seed[2198],seed[3725],seed[82],seed[1481],seed[7],seed[2629],seed[3033],seed[2019],seed[1507],seed[3184],seed[1885],seed[3354],seed[503],seed[2314],seed[3528],seed[1794],seed[3625],seed[4069],seed[3230],seed[3656],seed[704],seed[2533],seed[2476],seed[1399],seed[582],seed[1921],seed[3012],seed[976],seed[2768],seed[1831],seed[546],seed[3116],seed[4],seed[2468],seed[2056],seed[3325],seed[2095],seed[2154],seed[2396],seed[318],seed[270],seed[1007],seed[2559],seed[2924],seed[2706],seed[1477],seed[2998],seed[1945],seed[3010],seed[3066],seed[129],seed[2862],seed[3305],seed[722],seed[1423],seed[3319],seed[1879],seed[2292],seed[2547],seed[3142],seed[1968],seed[2508],seed[1754],seed[1607],seed[3879],seed[864],seed[1009],seed[2073],seed[417],seed[1636],seed[154],seed[2405],seed[2360],seed[3086],seed[2442],seed[3834],seed[2523],seed[1578],seed[148],seed[1107],seed[4047],seed[2756],seed[1491],seed[2558],seed[3810],seed[3568],seed[2981],seed[1790],seed[2970],seed[2366],seed[3576],seed[3799],seed[3893],seed[3600],seed[3803],seed[1245],seed[1461],seed[1005],seed[3418],seed[1054],seed[1194],seed[563],seed[765],seed[2192],seed[926],seed[2289],seed[1307],seed[1302],seed[3125],seed[289],seed[2929],seed[858],seed[3765],seed[3781],seed[806],seed[1235],seed[1695],seed[3490],seed[3398],seed[446],seed[1567],seed[1742],seed[1415],seed[299],seed[1716],seed[264],seed[538],seed[3875],seed[2514],seed[2015],seed[800],seed[3009],seed[3165],seed[1667],seed[2719],seed[2063],seed[398],seed[1411],seed[119],seed[4093],seed[2906],seed[2000],seed[3119],seed[643],seed[2661],seed[459],seed[1673],seed[3683],seed[1021],seed[3903],seed[1316],seed[3381],seed[527],seed[769],seed[2740],seed[3494],seed[1779],seed[2288],seed[1229],seed[2266],seed[995],seed[853],seed[1439],seed[3286],seed[4080],seed[3368],seed[334],seed[2807],seed[767],seed[3355],seed[77],seed[461],seed[949],seed[1963],seed[3429],seed[2551],seed[1941],seed[3155],seed[1125],seed[3178],seed[3107],seed[1455],seed[3570],seed[2861],seed[3995],seed[1610],seed[2042],seed[115],seed[2465],seed[179],seed[1803],seed[2787],seed[2565],seed[1094],seed[702],seed[2753],seed[3592],seed[287],seed[3851],seed[1694],seed[2087],seed[877],seed[1799],seed[3382],seed[1976],seed[3002],seed[258],seed[3708],seed[3272],seed[637],seed[2471],seed[3124],seed[1730],seed[2635],seed[3036],seed[513],seed[1661],seed[3684],seed[1375],seed[3709],seed[3587],seed[2168],seed[1185],seed[180],seed[197],seed[912],seed[76],seed[2299],seed[9],seed[683],seed[3136],seed[1015],seed[2698],seed[2483],seed[3615],seed[2026],seed[184],seed[1867],seed[1940],seed[2004],seed[132],seed[2274],seed[2053],seed[2572],seed[979],seed[1419],seed[843],seed[1624],seed[511],seed[3724],seed[68],seed[1269],seed[2995],seed[2790],seed[4009],seed[2939],seed[3548],seed[2632],seed[3941],seed[3222],seed[1965],seed[2333],seed[510],seed[176],seed[92],seed[2567],seed[4090],seed[3174],seed[711],seed[761],seed[768],seed[692],seed[3830],seed[2153],seed[2744],seed[474],seed[3866],seed[1715],seed[1565],seed[1562],seed[656],seed[1360],seed[2363],seed[1937],seed[3177],seed[888],seed[3435],seed[2530],seed[1807],seed[2391],seed[697],seed[654],seed[1982],seed[1322],seed[441],seed[165],seed[3839],seed[3602],seed[522],seed[653],seed[1713],seed[239],seed[2690],seed[1118],seed[1179],seed[2487],seed[1773],seed[1035],seed[2838],seed[4014],seed[991],seed[2061],seed[3881],seed[3118],seed[297],seed[885],seed[2488],seed[3651],seed[1719],seed[567],seed[2329],seed[1145],seed[1299],seed[2420],seed[2842],seed[472],seed[3442],seed[3763],seed[3361],seed[1109],seed[2562],seed[2003],seed[2017],seed[1449],seed[2328],seed[4021],seed[1698],seed[49],seed[2963],seed[1232],seed[3426],seed[2846],seed[3000],seed[1309],seed[191],seed[2824],seed[2648],seed[1866],seed[2207],seed[15],seed[1219],seed[2074],seed[2474],seed[1398],seed[228],seed[3309],seed[1336],seed[2452],seed[3397],seed[2879],seed[3812],seed[465],seed[1708],seed[3198],seed[416],seed[809],seed[61],seed[2209],seed[3658],seed[3678],seed[2702],seed[4007],seed[439],seed[3721],seed[2892],seed[1001],seed[2705],seed[1255],seed[2169],seed[2826],seed[2933],seed[3115],seed[1057],seed[1527],seed[2603],seed[1528],seed[2585],seed[2175],seed[1961],seed[1476],seed[101],seed[682],seed[3945],seed[2365],seed[2241],seed[2215],seed[3930],seed[1345],seed[2542],seed[2043],seed[504],seed[1922],seed[1193],seed[242],seed[1253],seed[1133],seed[1207],seed[341],seed[1936],seed[491],seed[507],seed[2305],seed[55],seed[1506],seed[4062],seed[3662],seed[3395],seed[3538],seed[1577],seed[1680],seed[4052],seed[1237],seed[2390],seed[2949],seed[1850],seed[2261],seed[897],seed[3789],seed[2406],seed[2269],seed[665],seed[971],seed[2774],seed[731],seed[1457],seed[2917],seed[996],seed[3451],seed[244],seed[2186],seed[2258],seed[1409],seed[1166],seed[948],seed[2358],seed[2236],seed[4020],seed[3955],seed[804],seed[2755],seed[4089],seed[201],seed[63],seed[2039],seed[3046],seed[1271],seed[719],seed[1775],seed[727],seed[2357],seed[3275],seed[1814],seed[862],seed[2089],seed[3065],seed[89],seed[3915],seed[1615],seed[2013],seed[1923],seed[2084],seed[218],seed[79],seed[1024],seed[2173],seed[2537],seed[3530],seed[3705],seed[4037],seed[486],seed[251],seed[23],seed[3205],seed[338],seed[2271],seed[3847],seed[2541],seed[676],seed[1746],seed[2229],seed[2115],seed[1918],seed[899],seed[2600],seed[3689],seed[1689],seed[3883],seed[1972],seed[2163],seed[3515],seed[480],seed[3001],seed[1920],seed[1117],seed[2232],seed[2254],seed[1004],seed[2426],seed[425],seed[389],seed[3711],seed[2735],seed[2421],seed[1508],seed[1066],seed[500],seed[3983],seed[4058],seed[570],seed[3506],seed[3285],seed[2934],seed[710],seed[3947],seed[3111],seed[2262],seed[3399],seed[73],seed[1887],seed[421],seed[3473],seed[3220],seed[268],seed[1261],seed[1137],seed[1721],seed[37],seed[2776],seed[3394],seed[3200],seed[2142],seed[1282],seed[2703],seed[667],seed[1784],seed[1592],seed[640],seed[3642],seed[3956],seed[3345],seed[720],seed[535],seed[3385],seed[2102],seed[1167],seed[1260],seed[3687],seed[1357],seed[3137],seed[2513],seed[3087],seed[2227],seed[2823],seed[2372],seed[2896],seed[1048],seed[3777],seed[3208],seed[4060],seed[790],seed[453],seed[3234],seed[1433],seed[766],seed[2076],seed[3535],seed[569],seed[3785],seed[688],seed[1640],seed[624],seed[3551],seed[1218],seed[1365],seed[1385],seed[3589],seed[3189],seed[3186],seed[1300],seed[3620],seed[20],seed[108],seed[2709],seed[2088],seed[122],seed[855],seed[125],seed[319],seed[2880],seed[1556],seed[3874],seed[2172],seed[4043],seed[447],seed[3547],seed[2282],seed[1127],seed[1581],seed[2213],seed[261],seed[2238],seed[2034],seed[658],seed[1816],seed[3655],seed[21],seed[1173],seed[2691],seed[2230],seed[541],seed[3402],seed[1099],seed[3288],seed[2516],seed[162],seed[1128],seed[3102],seed[212],seed[1381],seed[3173],seed[2371],seed[3612],seed[1489],seed[1389],seed[1583],seed[2991],seed[3202],seed[327],seed[884],seed[686],seed[2322],seed[357],seed[2831],seed[1039],seed[1430],seed[962],seed[1435],seed[3149],seed[3013],seed[1828],seed[3987],seed[3421],seed[3408],seed[3761],seed[3074],seed[3023],seed[3018],seed[3059],seed[3168],seed[568],seed[3140],seed[3801],seed[3112],seed[284],seed[1200],seed[2078],seed[2475],seed[2802],seed[88],seed[3984],seed[3105],seed[875],seed[1505],seed[3778],seed[785],seed[2313],seed[3386],seed[817],seed[2693],seed[2555],seed[1276],seed[2704],seed[4006],seed[1745],seed[243],seed[385],seed[2873],seed[810],seed[771],seed[2742],seed[966],seed[1956],seed[345],seed[3431],seed[2816],seed[2461],seed[1584],seed[3364],seed[1258],seed[1717],seed[3730],seed[1362],seed[1970],seed[1392],seed[198],seed[2440],seed[2489],seed[1871],seed[3281],seed[3324],seed[1536],seed[3921],seed[3938],seed[3206],seed[2291],seed[231],seed[3745],seed[3635],seed[178],seed[3121],seed[1198],seed[2504],seed[4071],seed[3608],seed[2145],seed[2553],seed[1888],seed[1662],seed[652],seed[1523],seed[1177],seed[3905],seed[4045],seed[104],seed[3850],seed[2161],seed[2875],seed[2779],seed[3936],seed[1599],seed[798],seed[2659],seed[661],seed[2660],seed[3719],seed[2930],seed[1537],seed[1981],seed[3299],seed[670],seed[2611],seed[2344],seed[1532],seed[2409],seed[2395],seed[2410],seed[350],seed[3567],seed[714],seed[3546],seed[707],seed[3466],seed[151],seed[2671],seed[2878],seed[410],seed[1143],seed[3317],seed[3741],seed[3271],seed[560],seed[1171],seed[1551],seed[2138],seed[3920],seed[2786],seed[65],seed[915],seed[826],seed[2552],seed[577],seed[3024],seed[2281],seed[3160],seed[2699],seed[2893],seed[1554],seed[3161],seed[3212],seed[247],seed[2350],seed[1418],seed[1056],seed[1600],seed[3563],seed[1726],seed[1657],seed[4079],seed[146],seed[2573],seed[2362],seed[3504],seed[2683],seed[3242],seed[2864],seed[1826],seed[3480],seed[2808],seed[3775],seed[1488],seed[3605],seed[2310],seed[3864],seed[3092],seed[3123],seed[870],seed[3353],seed[133],seed[2066],seed[2718],seed[748],seed[2948],seed[876],seed[1482],seed[1326],seed[3327],seed[337],seed[3463],seed[3910],seed[2979],seed[3918],seed[2710],seed[802],seed[2890],seed[3007],seed[1484],seed[657],seed[1652],seed[1518],seed[1631],seed[1856],seed[3562],seed[1511],seed[3372],seed[3210],seed[3630],seed[1767],seed[517],seed[3039],seed[1184],seed[646],seed[3641],seed[2940],seed[2863],seed[381],seed[1743],seed[130],seed[1142],seed[2277],seed[1350],seed[600],seed[1855],seed[46],seed[1055],seed[1804],seed[1479],seed[1911],seed[4040],seed[584],seed[255],seed[916],seed[3071],seed[689],seed[2459],seed[2195],seed[1722],seed[860],seed[782],seed[832],seed[1705],seed[3122],seed[3377],seed[1660],seed[537],seed[1327],seed[3088],seed[3986],seed[3307],seed[2759],seed[1230],seed[1646],seed[2577],seed[1215],seed[3289],seed[4082],seed[2877],seed[1601],seed[913],seed[3970],seed[2525],seed[3681],seed[2339],seed[2785],seed[3806],seed[3784],seed[1338],seed[846],seed[4027],seed[3179],seed[2761],seed[141],seed[3460],seed[1164],seed[1520],seed[3196],seed[2435],seed[323],seed[293],seed[2952],seed[2048],seed[87],seed[881],seed[3323],seed[3581],seed[762],seed[3979],seed[206],seed[3089],seed[2206],seed[3552],seed[458],seed[2033],seed[60],seed[1306],seed[2701],seed[2805],seed[155],seed[3972],seed[2545],seed[1513],seed[3467],seed[1312],seed[2355],seed[3751],seed[2256],seed[1901],seed[3294],seed[2912],seed[210],seed[2352],seed[585],seed[4070],seed[1546],seed[3326],seed[3128],seed[1793],seed[2598],seed[1603],seed[2393],seed[2347],seed[1737],seed[698],seed[3855],seed[3359],seed[1549],seed[428],seed[161],seed[1820],seed[558],seed[1622],seed[673],seed[2568],seed[1678],seed[3601],seed[1979],seed[1394],seed[1003],seed[2766],seed[669],seed[2308],seed[1633],seed[1666],seed[2092],seed[2490],seed[2343],seed[110],seed[3465],seed[1217],seed[71],seed[2472],seed[252],seed[2985],seed[1380],seed[588],seed[3621],seed[4054],seed[2609],seed[553],seed[2665],seed[2251],seed[1574],seed[200],seed[1458],seed[3176],seed[1079],seed[4064],seed[2764],seed[820],seed[2670],seed[887],seed[1440],seed[2085],seed[2788],seed[3080],seed[2211],seed[3097],seed[2664],seed[3491],seed[1865],seed[1621],seed[2607],seed[177],seed[1273],seed[118],seed[1720],seed[3900],seed[2116],seed[62],seed[1944],seed[1672],seed[573],seed[3130],seed[3223],seed[2590],seed[2321],seed[758],seed[1356],seed[1905],seed[2259],seed[3110],seed[2099],seed[3848],seed[3791],seed[935],seed[1490],seed[2159],seed[1036],seed[1061],seed[409],seed[2283],seed[796],seed[4087],seed[3943],seed[1420],seed[3558],seed[1605],seed[2300],seed[3297],seed[2891],seed[2216],seed[2515],seed[2280],seed[965],seed[1174],seed[1501],seed[550],seed[921],seed[911],seed[540],seed[375],seed[2898],seed[2369],seed[215],seed[1924],seed[625],seed[3019],seed[3409],seed[2141],seed[928],seed[2597],seed[2535],seed[460],seed[1596],seed[988],seed[3075],seed[2035],seed[3016],seed[647],seed[3557],seed[2257],seed[4013],seed[2849],seed[3419],seed[1031],seed[1303],seed[1050],seed[149],seed[3371],seed[1119],seed[111],seed[74],seed[2151],seed[1530],seed[3135],seed[3633],seed[3070],seed[156],seed[2639],seed[2682],seed[1453],seed[2713],seed[1759],seed[4072],seed[232],seed[4074],seed[3606],seed[2336],seed[38],seed[752],seed[2579],seed[1144],seed[1251],seed[1126],seed[2093],seed[2625],seed[3352],seed[1264],seed[2165],seed[3422],seed[2947],seed[3758],seed[325],seed[2070],seed[3675],seed[3591],seed[4050],seed[2375],seed[2136],seed[2593],seed[778],seed[1367],seed[986],seed[1279],seed[1747],seed[97],seed[3772],seed[3424],seed[3964],seed[246],seed[2543],seed[2315],seed[3704],seed[2117],seed[1585],seed[54],seed[2325],seed[424],seed[2255],seed[920],seed[361],seed[2578],seed[207],seed[2249],seed[4049],seed[3703],seed[2001],seed[128],seed[1116],seed[2411],seed[145],seed[506],seed[1785],seed[2407],seed[3583],seed[3807],seed[356],seed[2217],seed[1782],seed[3388],seed[775],seed[26],seed[592],seed[1899],seed[2673],seed[1211],seed[2994],seed[2874],seed[3996],seed[1731],seed[2399],seed[47],seed[304],seed[2902],seed[1542],seed[2707],seed[2630],seed[3434],seed[3503],seed[3197],seed[3030],seed[1620],seed[2131],seed[593],seed[3350],seed[1684],seed[3688],seed[992],seed[1602],seed[1131],seed[2587],seed[2750],seed[2794],seed[2678],seed[4035],seed[2905],seed[3497],seed[40],seed[3185],seed[2645],seed[1],seed[1157],seed[3259],seed[3433],seed[891],seed[2649],seed[3928],seed[3796],seed[3670],seed[2996],seed[565],seed[2058],seed[1777],seed[159],seed[2105],seed[3157],seed[2064],seed[1278],seed[777],seed[2278],seed[3269],seed[93],seed[2834],seed[2637],seed[937],seed[3407],seed[3489],seed[3525],seed[856],seed[2201],seed[2804],seed[1058],seed[2389],seed[3084],seed[534],seed[2051],seed[923],seed[2638],seed[2622],seed[1783],seed[1832],seed[1456],seed[2183],seed[1448],seed[1791],seed[1081],seed[3150],seed[548],seed[479],seed[2960],seed[1579],seed[1014],seed[351],seed[581],seed[1475],seed[1880],seed[3818],seed[4030],seed[1751],seed[476],seed[980],seed[3518],seed[1387],seed[1104],seed[2833],seed[1686],seed[1006],seed[3911],seed[3449],seed[1197],seed[332],seed[3493],seed[2810],seed[1796],seed[3573],seed[3985],seed[615],seed[1135],seed[2481],seed[2550],seed[3499],seed[743],seed[3366],seed[502],seed[2915],seed[1159],seed[1372],seed[1538],seed[418],seed[2049],seed[2723],seed[3582],seed[2443],seed[2770],seed[139],seed[2382],seed[2655],seed[2851],seed[85],seed[3935],seed[3586],seed[3152],seed[2999],seed[3896],seed[611],seed[2644],seed[3901],seed[2869],seed[2120],seed[2140],seed[1853],seed[2268],seed[3584],seed[613],seed[1960],seed[330],seed[1053],seed[42],seed[182],seed[1034],seed[1347],seed[2926],seed[2741],seed[505],seed[3646],seed[94],seed[2147],seed[773],seed[1216],seed[2446],seed[3697],seed[1894],seed[2096],seed[2936],seed[2643],seed[716],seed[137],seed[982],seed[2867],seed[2414],seed[865],seed[377],seed[2046],seed[328],seed[572],seed[1366],seed[3108],seed[1861],seed[1335],seed[2265],seed[2646],seed[2956],seed[533],seed[3191],seed[1374],seed[1948],seed[3731],seed[285],seed[1246],seed[3256],seed[2663],seed[3578],seed[1971],seed[750],seed[2006],seed[3254],seed[164],seed[436],seed[1844],seed[3332],seed[1916],seed[784],seed[3120],seed[1331],seed[397],seed[898],seed[3396],seed[852],seed[2495],seed[172],seed[371],seed[3968],seed[2941],seed[2028],seed[1065],seed[2641],seed[3695],seed[1572],seed[1890],seed[29],seed[170],seed[622],seed[1644],seed[954],seed[2528],seed[1120],seed[1692],seed[1874],seed[2221],seed[2858],seed[3529],seed[1813],seed[1738],seed[4055],seed[2773],seed[3203],seed[833],seed[934],seed[4023],seed[770],seed[1780],seed[2675],seed[612],seed[2604],seed[158],seed[1909],seed[1649],seed[3767],seed[759],seed[2983],seed[2243],seed[1575],seed[1016],seed[854],seed[3038],seed[751],seed[2927],seed[1727],seed[3669],seed[999],seed[2584],seed[3311],seed[3991],seed[217],seed[114],seed[3835],seed[3842],seed[3117],seed[1829],seed[2922],seed[3759],seed[1707],seed[873],seed[2463],seed[1115],seed[1139],seed[2818],seed[1550],seed[3443],seed[3824],seed[2456],seed[1852],seed[4084],seed[3474],seed[4008],seed[1140],seed[1002],seed[3664],seed[1709],seed[1823],seed[890],seed[946],seed[649],seed[2497],seed[124],seed[2129],seed[3415],seed[1351],seed[1632],seed[1228],seed[2137],seed[3049],seed[3942],seed[1369],seed[402],seed[3427],seed[2582],seed[3723],seed[390],seed[223],seed[1630],seed[3069],seed[3461],seed[1122],seed[3251],seed[3944],seed[2174],seed[2510],seed[1926],seed[369],seed[443],seed[3701],seed[2606],seed[2245],seed[2155],seed[3769],seed[1953],seed[2478],seed[3237],seed[863],seed[1358],seed[2052],seed[3280],seed[3965],seed[1676],seed[717],seed[2021],seed[3571],seed[1869],seed[3329],seed[2381],seed[1744],seed[3008],seed[1098],seed[3126],seed[942],seed[2684],seed[3405],seed[3509],seed[406],seed[1992],seed[559],seed[2397],seed[478],seed[3904],seed[1540],seed[2285],seed[163],seed[3783],seed[774],seed[3978],seed[1494],seed[1771],seed[2486],seed[3260],seed[3960],seed[157],seed[1900],seed[3005],seed[2975],seed[423],seed[970],seed[1121],seed[1332],seed[358],seed[3829],seed[3502],seed[1170],seed[744],seed[3610],seed[2509],seed[849],seed[2128],seed[857],seed[83],seed[981],seed[664],seed[1041],seed[1723],seed[1974],seed[320],seed[1202],seed[2812],seed[578],seed[471],seed[3238],seed[3629],seed[2246],seed[1408],seed[3423],seed[932],seed[2342],seed[2965],seed[1765],seed[1576],seed[3981],seed[1262],seed[1841],seed[1199],seed[963],seed[2388],seed[1178],seed[2666],seed[2796],seed[2210],seed[1247],seed[3457],seed[1623],seed[3523],seed[3786],seed[3127],seed[772],seed[691],seed[2799],seed[2466],seed[3828],seed[1405],seed[1802],seed[395],seed[99],seed[690],seed[2712],seed[2653],seed[2367],seed[455],seed[1589],seed[1864],seed[958],seed[2149],seed[1642],seed[1499],seed[997],seed[3585],seed[3390],seed[1996],seed[3143],seed[2913],seed[4017],seed[3148],seed[2844],seed[1792],seed[3363],seed[1183],seed[2467],seed[194],seed[2214],seed[3753],seed[3845],seed[1428],seed[3468],seed[1180],seed[1010],seed[3926],seed[1821],seed[2674],seed[70],seed[3109],seed[2942],seed[1653],seed[3296],seed[626],seed[1770],seed[1298],seed[2260],seed[1973],seed[2044],seed[3091],seed[726],seed[1984],seed[1187],seed[2687],seed[2177],seed[2018],seed[2726],seed[2730],seed[2082],seed[3543],seed[2250],seed[1346],seed[309],seed[238],seed[2364],seed[3762],seed[2445],seed[1704],seed[3887],seed[894],seed[493],seed[3980],seed[1132],seed[3351],seed[1516],seed[2432],seed[4092],seed[2914],seed[3063],seed[3510],seed[1641],seed[374],seed[909],seed[143],seed[2077],seed[2885],seed[2020],seed[3660],seed[3726],seed[3282],seed[824],seed[2919],seed[1256],seed[3954],seed[2057],seed[2524],seed[28],seed[3609],seed[1325],seed[2002],seed[3884],seed[1487],seed[1854],seed[3895],seed[2112],seed[2784],seed[2431],seed[1496],seed[2668],seed[3802],seed[2007],seed[1849],seed[2040],seed[2506],seed[1123],seed[3146],seed[524],seed[2309],seed[1165],seed[1733],seed[757],seed[51],seed[2132],seed[2290],seed[80],seed[3952],seed[604],seed[952],seed[3872],seed[2114],seed[3973],seed[3414],seed[1000],seed[3545],seed[2180],seed[866],seed[3513],seed[536],seed[3225],seed[1480],seed[3702],seed[3483],seed[1434],seed[552],seed[4036],seed[1227],seed[4073],seed[1568],seed[3686],seed[1729],seed[2647],seed[213],seed[3556],seed[462],seed[2688],seed[1275],seed[1701],seed[556],seed[2143],seed[3696],seed[383],seed[3077],seed[2957],seed[3204],seed[677],seed[1426],seed[606],seed[8],seed[848],seed[4005],seed[1402],seed[1416],seed[2560],seed[1208],seed[614],seed[3857],seed[32],seed[2331],seed[1314],seed[1321],seed[1580],seed[3195],seed[2403],seed[3247],seed[3682],seed[274],seed[4086],seed[3035],seed[674],seed[3060],seed[401],seed[3261],seed[1500],seed[2962],seed[2621],seed[1444],seed[1495],seed[3101],seed[2782],seed[1582],seed[3690],seed[1502],seed[3383],seed[407],seed[1711],seed[1076],seed[2303],seed[709],seed[3707],seed[98],seed[127],seed[382],seed[1553],seed[1761],seed[2394],seed[2809],seed[5],seed[3134],seed[2566],seed[3347],seed[2832],seed[2197],seed[3450],seed[3746],seed[1818],seed[3680],seed[2840],seed[1284],seed[1836],seed[3643],seed[2450],seed[1725],seed[1519],seed[3293],seed[2424],seed[708],seed[984],seed[1288],seed[1364],seed[3058],seed[3950],seed[1101],seed[354],seed[1685],seed[3335],seed[2376],seed[189],seed[3892],seed[22],seed[3880],seed[2184],seed[4057],seed[699],seed[2247],seed[3213],seed[497],seed[601],seed[922],seed[3430],seed[1295],seed[2897],seed[66],seed[1267],seed[3055],seed[2242],seed[3428],seed[1146],seed[109],seed[1617],seed[2298],seed[286],seed[3050],seed[1152],seed[1668],seed[1859],seed[336],seed[2098],seed[3479],seed[3663],seed[695],seed[2359],seed[3444],seed[2301],seed[1712],seed[1445],seed[451],seed[185],seed[718],seed[2751],seed[431],seed[3631],seed[3246],seed[3649],seed[1564],seed[1195],seed[3056],seed[896],seed[2423],seed[3215],seed[147],seed[91],seed[2297],seed[3840],seed[1503],seed[3899],seed[3932],seed[840],seed[2697],seed[2152],seed[426],seed[1393],seed[2430],seed[4010],seed[3257],seed[1635],seed[380],seed[31],seed[367],seed[2904],seed[3738],seed[780],seed[1379],seed[353],seed[1096],seed[3712],seed[3072],seed[187],seed[64],seed[1220],seed[2279],seed[3478],seed[3760],seed[2133],seed[2669],seed[1654],seed[1090],seed[2496],seed[783],seed[1703],seed[3106],seed[3644],seed[1959],seed[1340],seed[2589],seed[3315],seed[1371],seed[2617],seed[2224],seed[3774],seed[314],seed[776],seed[532],seed[276],seed[494],seed[3253],seed[2103],seed[241],seed[3241],seed[1138],seed[1786],seed[1293],seed[3201],seed[631],seed[250],seed[2888],seed[1105],seed[1656],seed[1033],seed[1758],seed[2819],seed[1388],seed[144],seed[740],seed[2856],seed[1958],seed[1071],seed[960],seed[2387],seed[2850],seed[3331],seed[1051],seed[3373],seed[2008],seed[2841],seed[365],seed[3517],seed[3750],seed[1679],seed[52],seed[1319],seed[399],seed[3797],seed[2437],seed[19],seed[1919],seed[457],seed[910],seed[967],seed[271],seed[2032],seed[2767],seed[1691],seed[1877],seed[482],seed[1964],seed[1311],seed[1999],seed[823],seed[2055],seed[4024],seed[1280],seed[2583],seed[2845],seed[555],seed[666],seed[3263],seed[86],seed[2814],seed[3219],seed[3511],seed[3953],seed[760],seed[610],seed[1993],seed[279],seed[3626],seed[414],seed[3624],seed[3961],seed[2449],seed[3476],seed[100],seed[3015],seed[468],seed[721],seed[2988],seed[1728],seed[2222],seed[737],seed[3349],seed[514],seed[3477],seed[1892],seed[2187],seed[1862],seed[3815],seed[0],seed[2576],seed[2791],seed[1891],seed[90],seed[2827],seed[1498],seed[4039],seed[168],seed[1591],seed[847],seed[3472],seed[2494],seed[930],seed[3833],seed[2758],seed[419],seed[2124],seed[630],seed[1286],seed[1983],seed[2716],seed[1619],seed[1296],seed[3539],seed[3794],seed[703],seed[3095],seed[2083],seed[2402],seed[1812],seed[1990],seed[2263],seed[1706],seed[1955],seed[1422],seed[3226],seed[2160],seed[501],seed[134],seed[321],seed[17],seed[3598],seed[1093],seed[3971],seed[387],seed[1270],seed[1535],seed[3982],seed[3365],seed[2239],seed[2997],seed[822],seed[496],seed[1967],seed[2024],seed[3969],seed[723],seed[907],seed[3648],seed[290],seed[2657],seed[2068],seed[3268],seed[4044],seed[263],seed[1756],seed[745],seed[1473],seed[2538],seed[1566],seed[2591],seed[2200],seed[1470],seed[1655],seed[2775],seed[275],seed[3236],seed[413],seed[2859],seed[490],seed[2094],seed[3054],seed[126],seed[442],seed[786],seed[1329],seed[1224],seed[2554],seed[3240],seed[2640],seed[2821],seed[1072],seed[1181],seed[1886],seed[819],seed[1466],seed[2752],seed[1534],seed[3958],seed[2564],seed[2870],seed[57],seed[3674],seed[2757],seed[2059],seed[3166],seed[4032],seed[214],seed[869],seed[1318],seed[861],seed[2171],seed[2866],seed[781],seed[587],seed[1932],seed[1469],seed[940],seed[292],seed[2521],seed[3369],seed[730],seed[1618],seed[498],seed[3042],seed[3531],seed[1337],seed[2793],seed[282],seed[3132],seed[3507],seed[2626],seed[3052],seed[2451],seed[1027],seed[3808],seed[4012],seed[3940],seed[1734],seed[2580],seed[3617],seed[3180],seed[386],seed[1313],seed[4083],seed[2134],seed[342],seed[3715],seed[1805],seed[388],seed[470],seed[192],seed[363],seed[3448],seed[1080],seed[1342],seed[1732],seed[2100],seed[234],seed[1969],seed[2769],seed[2248],seed[1088],seed[641],seed[2938],seed[3865],seed[1858],seed[1989],seed[1611],seed[3182],seed[2030],seed[1410],seed[1609],seed[3459],seed[1100],seed[2419],seed[1837],seed[1196],seed[1268],seed[3650],seed[2418],seed[671],seed[3768],seed[3838],seed[2571],seed[3047],seed[1659],seed[2188],seed[1638],seed[825],seed[3078],seed[1413],seed[2815],seed[3412],seed[1724],seed[2781],seed[450],seed[2493],seed[554],seed[2434],seed[2284],seed[3290],seed[1898],seed[1169],seed[1896],seed[2534],seed[3819],seed[3048],seed[379],seed[3754],seed[2144],seed[3885],seed[3156],seed[1162],seed[1760],seed[3638],seed[3011],seed[3685],seed[2462],seed[3114],seed[974],seed[340],seed[3057],seed[3856],seed[1020],seed[3262],seed[1062],seed[2353],seed[794],seed[2025],seed[1158],seed[3988],seed[1639],seed[2237],seed[1287],seed[2079],seed[226],seed[639],seed[2016],seed[3622],seed[3949],seed[1977],seed[1808],seed[3447],seed[4025],seed[1778],seed[2800],seed[2205],seed[1810],seed[3919],seed[1148],seed[2108],seed[1429],seed[2060],seed[2955],seed[2772],seed[1914],seed[1893],seed[3342],seed[3235],seed[3722],seed[2642],seed[1240],seed[1822],seed[245],seed[938],seed[994],seed[2212],seed[2920],seed[3618],seed[635],seed[1927],seed[713],seed[3340],seed[3853],seed[2304],seed[2398],seed[3163],seed[3028],seed[1710],seed[3521],seed[2199],seed[2065],seed[2307],seed[169],seed[3227],seed[3923],seed[1354],seed[3718],seed[3044],seed[1176],seed[4038],seed[1334],seed[2634],seed[464],seed[3889],seed[2724],seed[3099],seed[3244],seed[3728],seed[1878],seed[225],seed[1840],seed[3252],seed[596],seed[4031],seed[2820],seed[2803],seed[1212],seed[2620],seed[1857],seed[3094],seed[2233],seed[729],seed[310],seed[1441],seed[135],seed[487],seed[3471],seed[3239],seed[56],seed[4081],seed[348],seed[2253],seed[3813],seed[2903],seed[959],seed[3671],seed[1464],seed[2139],seed[874],seed[2416],seed[4042],seed[1570],seed[2778],seed[903],seed[6],seed[492],seed[1497],seed[2725],seed[914],seed[2749],seed[3387],seed[944],seed[2540],seed[333],seed[2931],seed[3634],seed[839],seed[1755],seed[2377],seed[1149],seed[2511],seed[186],seed[3579],seed[1616],seed[828],seed[3270],seed[3248],seed[638],seed[3541],seed[2320],seed[229],seed[195],seed[2966],seed[838],seed[4000],seed[3064],seed[3793],seed[235],seed[3188],seed[3732],seed[366],seed[3549],seed[2235],seed[3854],seed[50],seed[2429],seed[3481],seed[3512],seed[983],seed[2624],seed[483],seed[433],seed[2491],seed[1693],seed[437],seed[2146],seed[1817],seed[648],seed[3522],seed[3770],seed[3154],seed[4091],seed[2482],seed[3959],seed[3308],seed[1951],seed[508],seed[927],seed[700],seed[2715],seed[2127],seed[2876],seed[574],seed[2485],seed[632],seed[545],seed[3169],seed[3520],seed[893],seed[1669],seed[801],seed[485],seed[378],seed[2546],seed[1407],seed[668],seed[608],seed[3314],seed[495],seed[1204],seed[2386],seed[3998],seed[2680],seed[3131],seed[589],seed[3043],seed[1748],seed[3679],seed[3183],seed[1845],seed[2569],seed[3141],seed[3614],seed[2518],seed[889],seed[2507],seed[3604],seed[3344],seed[2413],seed[2522],seed[2570],seed[3897],seed[3809],seed[1089],seed[3749],seed[224],seed[3966],seed[808],seed[400],seed[3596],seed[3300],seed[368],seed[1904],seed[2351],seed[3826],seed[1827],seed[1903],seed[1403],seed[2935],seed[2992],seed[2631],seed[449],seed[1203],seed[1682],seed[2010],seed[2696],seed[3735],seed[2722],seed[2422],seed[998],seed[3594],seed[3729],seed[1236],seed[969],seed[1086],seed[4051],seed[3190],seed[1627],seed[842],seed[939],seed[3667],seed[2720],seed[850],seed[595],seed[2601],seed[3565],seed[1052],seed[872],seed[2505],seed[696],seed[3266],seed[705],seed[1028],seed[2041],seed[2519],seed[1571],seed[1994],seed[3167],seed[679],seed[2317],seed[4026],seed[2946],seed[2909],seed[2717],seed[3743],seed[3004],seed[3287],seed[1324],seed[3193],seed[598],seed[1047],seed[3475],seed[1848],seed[918],seed[724],seed[3367],seed[3455],seed[2189],seed[3488],seed[924],seed[2385],seed[1811],seed[2605],seed[183],seed[2792],seed[2974],seed[430],seed[2672],seed[1214],seed[3640],seed[583],seed[3836],seed[1084],seed[3569],seed[1222],seed[2130],seed[931],seed[1493],seed[3337],seed[2080],seed[272],seed[2900],seed[3909],seed[4095],seed[2374],seed[1868],seed[349],seed[204],seed[160],seed[2498],seed[2427],seed[3375],seed[3250],seed[257],seed[2839],seed[1555],seed[978],seed[3871],seed[355],seed[1182],seed[3931],seed[488],seed[3860],seed[1438],seed[1301],seed[557],seed[3665],seed[106],seed[1097],seed[1472],seed[807],seed[295],seed[254],seed[335],seed[3199],seed[2480],seed[2695],seed[445],seed[1797],seed[3380],seed[1658],seed[3221],seed[2327],seed[1384],seed[2323],seed[4094],seed[687],seed[3341],seed[3906],seed[259],seed[964],seed[1514],seed[3559],seed[2958],seed[1541],seed[2223],seed[2588],seed[3277],seed[693],seed[2685],seed[756],seed[3908],seed[818],seed[1044],seed[2731],seed[2106],seed[3139],seed[3554],seed[797],seed[3192],seed[4041],seed[1075],seed[835],seed[2737],seed[1986],seed[2031],seed[1414],seed[1544],seed[203],seed[2417],seed[3283],seed[3482],seed[1586],seed[3800],seed[3312],seed[1064],seed[1290],seed[3318],seed[663],seed[3073],seed[1690],seed[3771],seed[393],seed[3977],seed[2943],seed[3313],seed[779],seed[2536],seed[2150],seed[24],seed[3555],seed[404],seed[878],seed[4016],seed[3790],seed[2557],seed[2734],seed[1112],seed[3170],seed[405],seed[3795],seed[3623],seed[3566],seed[2477],seed[1025],seed[3310],seed[1697],seed[1370],seed[1073],seed[1460],seed[2341],seed[2464],seed[1884],seed[3844],seed[2473],seed[2368],seed[1947],seed[3742],seed[1049],seed[1315],seed[1085],seed[199],seed[516],seed[1650],seed[1504],seed[2881],seed[755],seed[3362],seed[3322],seed[1323],seed[586],seed[2244],seed[3438],seed[3659],seed[956],seed[2428],seed[269],seed[901],seed[3994],seed[1383],seed[2126],seed[3181],seed[1766],seed[3876],seed[3992],seed[1991],seed[3391],seed[2733],seed[1153],seed[1134],seed[2837],seed[2855],seed[2062],seed[152],seed[1946],seed[950],seed[448],seed[1424],seed[3948],seed[2780],seed[3229],seed[2899],seed[3744],seed[2918]}),
        .cross_prob(cross_prob),
        .codeword(codeword5),
        .received(received5)
        );
    
    bsc bsc6(
        .clk(clk),
        .reset(reset),
        .seed({seed[3333],seed[1882],seed[2180],seed[1478],seed[347],seed[3824],seed[9],seed[1363],seed[1908],seed[2134],seed[2917],seed[2601],seed[4038],seed[2948],seed[3576],seed[2516],seed[3599],seed[1370],seed[1913],seed[1089],seed[3313],seed[1462],seed[2216],seed[492],seed[1912],seed[1024],seed[3045],seed[3510],seed[909],seed[252],seed[3377],seed[3179],seed[587],seed[1482],seed[1396],seed[1835],seed[1866],seed[1997],seed[1278],seed[2660],seed[2382],seed[851],seed[3964],seed[1839],seed[2447],seed[2776],seed[864],seed[3194],seed[680],seed[359],seed[613],seed[1410],seed[1124],seed[2529],seed[2806],seed[3679],seed[3043],seed[519],seed[2589],seed[2804],seed[4050],seed[1394],seed[1144],seed[161],seed[125],seed[767],seed[3307],seed[4082],seed[2977],seed[2003],seed[3253],seed[4077],seed[3471],seed[3230],seed[3488],seed[154],seed[2843],seed[3072],seed[1443],seed[3055],seed[1461],seed[1915],seed[1353],seed[1250],seed[1006],seed[2118],seed[3139],seed[2068],seed[1776],seed[1179],seed[4063],seed[3823],seed[1760],seed[972],seed[391],seed[2527],seed[726],seed[228],seed[112],seed[245],seed[500],seed[1115],seed[3845],seed[581],seed[1890],seed[2803],seed[429],seed[2832],seed[2787],seed[870],seed[3787],seed[3640],seed[3722],seed[2188],seed[461],seed[2793],seed[1301],seed[2288],seed[2189],seed[2570],seed[3171],seed[2822],seed[3478],seed[3835],seed[3792],seed[298],seed[3019],seed[3553],seed[2362],seed[50],seed[3669],seed[1509],seed[3033],seed[1737],seed[1031],seed[1649],seed[3305],seed[3991],seed[1495],seed[1650],seed[2119],seed[771],seed[2884],seed[2503],seed[2786],seed[617],seed[3858],seed[1824],seed[1429],seed[596],seed[996],seed[46],seed[1576],seed[232],seed[559],seed[85],seed[974],seed[3592],seed[1075],seed[2468],seed[1718],seed[3147],seed[3632],seed[1813],seed[3736],seed[1193],seed[4040],seed[3409],seed[3235],seed[1800],seed[2761],seed[676],seed[1874],seed[3187],seed[1052],seed[2092],seed[1037],seed[3495],seed[1397],seed[2359],seed[631],seed[2102],seed[643],seed[2878],seed[4011],seed[2038],seed[3695],seed[3862],seed[2401],seed[2831],seed[1766],seed[714],seed[3976],seed[1785],seed[355],seed[3001],seed[2421],seed[1816],seed[1349],seed[250],seed[1273],seed[2735],seed[3412],seed[1811],seed[3830],seed[2290],seed[1696],seed[1621],seed[964],seed[3343],seed[1023],seed[2056],seed[1610],seed[3786],seed[1085],seed[2898],seed[2683],seed[2959],seed[603],seed[1653],seed[2133],seed[2823],seed[799],seed[3838],seed[2517],seed[3465],seed[3366],seed[3295],seed[3829],seed[3500],seed[2053],seed[3827],seed[2173],seed[2954],seed[947],seed[3924],seed[3586],seed[2870],seed[2961],seed[1065],seed[2137],seed[418],seed[442],seed[128],seed[313],seed[1463],seed[898],seed[1294],seed[412],seed[2398],seed[991],seed[1266],seed[1688],seed[2992],seed[755],seed[3116],seed[258],seed[805],seed[3330],seed[2923],seed[2391],seed[3997],seed[3698],seed[3107],seed[1487],seed[163],seed[1257],seed[2183],seed[1859],seed[143],seed[3565],seed[139],seed[1377],seed[3548],seed[3590],seed[1526],seed[748],seed[2984],seed[3987],seed[3185],seed[1472],seed[3563],seed[3146],seed[259],seed[620],seed[4062],seed[1086],seed[2711],seed[1585],seed[957],seed[2349],seed[1909],seed[1947],seed[2813],seed[3387],seed[2494],seed[2629],seed[2333],seed[2368],seed[2895],seed[2700],seed[3371],seed[3690],seed[1562],seed[990],seed[1427],seed[3524],seed[1697],seed[281],seed[80],seed[2544],seed[1107],seed[2689],seed[4078],seed[529],seed[1473],seed[2669],seed[1035],seed[3110],seed[1453],seed[1715],seed[2746],seed[4047],seed[200],seed[2591],seed[155],seed[1063],seed[3952],seed[1387],seed[1214],seed[3340],seed[1860],seed[3096],seed[448],seed[4018],seed[1351],seed[1002],seed[3130],seed[2040],seed[4004],seed[2723],seed[3948],seed[1659],seed[286],seed[2587],seed[89],seed[60],seed[2267],seed[1008],seed[1259],seed[3250],seed[826],seed[2082],seed[850],seed[2900],seed[215],seed[253],seed[729],seed[1579],seed[3483],seed[1440],seed[3456],seed[761],seed[1428],seed[1941],seed[1522],seed[815],seed[2017],seed[1898],seed[1442],seed[2208],seed[2159],seed[3814],seed[1729],seed[3803],seed[3405],seed[892],seed[396],seed[1983],seed[1437],seed[3419],seed[3125],seed[2609],seed[644],seed[1602],seed[1230],seed[3919],seed[1044],seed[1264],seed[3181],seed[3982],seed[763],seed[443],seed[690],seed[1403],seed[1594],seed[1596],seed[2511],seed[1080],seed[759],seed[2260],seed[2120],seed[3246],seed[509],seed[2552],seed[3438],seed[3353],seed[899],seed[1812],seed[3770],seed[160],seed[3003],seed[3937],seed[336],seed[3200],seed[710],seed[822],seed[2165],seed[3754],seed[1549],seed[692],seed[3023],seed[3008],seed[528],seed[829],seed[3011],seed[2280],seed[394],seed[2322],seed[2123],seed[1540],seed[4044],seed[2300],seed[1752],seed[3822],seed[1418],seed[3032],seed[3990],seed[2801],seed[756],seed[2231],seed[133],seed[3009],seed[3431],seed[873],seed[3121],seed[1064],seed[1553],seed[1498],seed[3082],seed[454],seed[1480],seed[2833],seed[126],seed[2073],seed[2840],seed[516],seed[1245],seed[2004],seed[3598],seed[1010],seed[2628],seed[356],seed[874],seed[1682],seed[3680],seed[3541],seed[3306],seed[1558],seed[1804],seed[769],seed[1846],seed[3931],seed[3463],seed[2987],seed[3207],seed[1185],seed[2905],seed[1571],seed[196],seed[293],seed[309],seed[1788],seed[1445],seed[730],seed[705],seed[2638],seed[1244],seed[1197],seed[3382],seed[2561],seed[1489],seed[2002],seed[1255],seed[1588],seed[518],seed[1077],seed[1676],seed[1960],seed[2268],seed[2950],seed[435],seed[1022],seed[181],seed[4056],seed[172],seed[2025],seed[3604],seed[3649],seed[3543],seed[3544],seed[3869],seed[3445],seed[3000],seed[1680],seed[3467],seed[1743],seed[101],seed[1105],seed[1793],seed[3605],seed[918],seed[876],seed[307],seed[3566],seed[2528],seed[2171],seed[2645],seed[2388],seed[2730],seed[1236],seed[917],seed[3837],seed[642],seed[928],seed[4070],seed[3358],seed[1864],seed[3167],seed[2373],seed[436],seed[3153],seed[4064],seed[800],seed[3221],seed[3715],seed[746],seed[1569],seed[3917],seed[2124],seed[2575],seed[3711],seed[1668],seed[2410],seed[3086],seed[510],seed[3391],seed[2579],seed[2569],seed[3112],seed[3567],seed[1829],seed[2886],seed[3572],seed[408],seed[602],seed[494],seed[2078],seed[2360],seed[2199],seed[3944],seed[3069],seed[2145],seed[1740],seed[2258],seed[2877],seed[2968],seed[1707],seed[3089],seed[1645],seed[3460],seed[929],seed[3458],seed[213],seed[2254],seed[741],seed[2089],seed[270],seed[3847],seed[2847],seed[3122],seed[579],seed[69],seed[3994],seed[1981],seed[2719],seed[2342],seed[3385],seed[1275],seed[2924],seed[859],seed[3354],seed[3036],seed[2475],seed[3658],seed[3998],seed[2224],seed[4080],seed[473],seed[27],seed[1239],seed[2734],seed[1441],seed[2936],seed[2939],seed[0],seed[66],seed[2705],seed[2146],seed[3664],seed[666],seed[3712],seed[2928],seed[1938],seed[2027],seed[3969],seed[2181],seed[3141],seed[2602],seed[2327],seed[831],seed[30],seed[3224],seed[824],seed[983],seed[1739],seed[624],seed[3346],seed[87],seed[1593],seed[3550],seed[1231],seed[238],seed[227],seed[1665],seed[3893],seed[3643],seed[2088],seed[2084],seed[1550],seed[2862],seed[2346],seed[1714],seed[306],seed[206],seed[2899],seed[1263],seed[2396],seed[1590],seed[3242],seed[3925],seed[205],seed[3015],seed[1510],seed[2670],seed[3891],seed[2577],seed[3562],seed[95],seed[959],seed[839],seed[3345],seed[3046],seed[1268],seed[4003],seed[1127],seed[37],seed[244],seed[1867],seed[3007],seed[3648],seed[361],seed[1606],seed[3192],seed[290],seed[1206],seed[2625],seed[1822],seed[1880],seed[1116],seed[2681],seed[424],seed[1184],seed[3198],seed[3904],seed[486],seed[2518],seed[3965],seed[989],seed[177],seed[3555],seed[1333],seed[267],seed[531],seed[593],seed[1644],seed[2110],seed[312],seed[1546],seed[444],seed[1012],seed[2174],seed[1056],seed[2011],seed[1651],seed[1156],seed[2458],seed[2469],seed[2428],seed[695],seed[628],seed[536],seed[4085],seed[760],seed[1026],seed[1166],seed[366],seed[954],seed[1987],seed[3499],seed[1485],seed[1152],seed[3859],seed[1280],seed[320],seed[662],seed[1066],seed[2452],seed[4072],seed[1316],seed[977],seed[1218],seed[2026],seed[3582],seed[1209],seed[1154],seed[2588],seed[4008],seed[610],seed[1533],seed[682],seed[1327],seed[1384],seed[1774],seed[2777],seed[465],seed[3962],seed[2942],seed[1420],seed[3947],seed[527],seed[470],seed[2805],seed[2467],seed[2827],seed[1270],seed[41],seed[1934],seed[3208],seed[3481],seed[23],seed[114],seed[3935],seed[1458],seed[1642],seed[2385],seed[2715],seed[1059],seed[2824],seed[2739],seed[265],seed[1452],seed[1771],seed[1222],seed[1667],seed[3867],seed[341],seed[3180],seed[2901],seed[49],seed[2604],seed[3621],seed[1552],seed[2999],seed[1286],seed[3915],seed[2855],seed[3812],seed[251],seed[2434],seed[4083],seed[3482],seed[3154],seed[226],seed[2741],seed[2355],seed[3772],seed[3178],seed[3031],seed[4052],seed[2210],seed[1974],seed[2639],seed[1019],seed[936],seed[2230],seed[131],seed[1221],seed[2616],seed[3341],seed[1271],seed[2631],seed[2808],seed[1272],seed[310],seed[1990],seed[2857],seed[728],seed[3685],seed[1732],seed[693],seed[285],seed[890],seed[2724],seed[2269],seed[2876],seed[2606],seed[2894],seed[3357],seed[3166],seed[3209],seed[2851],seed[81],seed[604],seed[1611],seed[3150],seed[168],seed[333],seed[3229],seed[330],seed[167],seed[1702],seed[3101],seed[1337],seed[3104],seed[3188],seed[493],seed[1910],seed[452],seed[2885],seed[194],seed[1305],seed[2546],seed[4071],seed[2433],seed[1207],seed[3049],seed[1111],seed[3367],seed[3558],seed[3068],seed[2212],seed[153],seed[3570],seed[2585],seed[655],seed[346],seed[1917],seed[2223],seed[938],seed[3175],seed[76],seed[2315],seed[3421],seed[2214],seed[411],seed[1252],seed[354],seed[3173],seed[1748],seed[3284],seed[506],seed[3352],seed[2324],seed[2654],seed[2913],seed[3725],seed[1946],seed[337],seed[2105],seed[1138],seed[2108],seed[2063],seed[3073],seed[1005],seed[875],seed[2242],seed[3578],seed[3677],seed[236],seed[209],seed[340],seed[2232],seed[539],seed[900],seed[2972],seed[637],seed[1499],seed[2736],seed[317],seed[3155],seed[2170],seed[3136],seed[2157],seed[462],seed[2249],seed[382],seed[1970],seed[284],seed[269],seed[1781],seed[3797],seed[1210],seed[3940],seed[1400],seed[2997],seed[1963],seed[1520],seed[2557],seed[2096],seed[3312],seed[2062],seed[2679],seed[3678],seed[2465],seed[4074],seed[2257],seed[667],seed[15],seed[3355],seed[1158],seed[3608],seed[525],seed[3767],seed[3035],seed[2168],seed[2023],seed[2309],seed[201],seed[2295],seed[1455],seed[1741],seed[2226],seed[2633],seed[272],seed[1574],seed[659],seed[2772],seed[2329],seed[843],seed[3241],seed[1148],seed[53],seed[1758],seed[2485],seed[722],seed[798],seed[220],seed[453],seed[1],seed[1889],seed[944],seed[379],seed[1556],seed[198],seed[397],seed[2526],seed[908],seed[3879],seed[3957],seed[2237],seed[2816],seed[63],seed[86],seed[3138],seed[1841],seed[552],seed[1627],seed[3328],seed[3084],seed[2201],seed[975],seed[3875],seed[2412],seed[1968],seed[846],seed[3557],seed[3067],seed[2731],seed[3260],seed[127],seed[3507],seed[1634],seed[2795],seed[2982],seed[542],seed[3574],seed[2826],seed[1362],seed[119],seed[3790],seed[1411],seed[1899],seed[4067],seed[491],seed[3734],seed[2944],seed[1046],seed[1000],seed[3403],seed[1117],seed[1773],seed[274],seed[2172],seed[2319],seed[2314],seed[3014],seed[2690],seed[554],seed[3968],seed[2983],seed[3849],seed[994],seed[952],seed[1720],seed[3381],seed[384],seed[3936],seed[1211],seed[387],seed[35],seed[2325],seed[3816],seed[499],seed[3317],seed[3102],seed[568],seed[2044],seed[16],seed[249],seed[428],seed[3047],seed[3581],seed[1421],seed[2219],seed[3441],seed[386],seed[1199],seed[3446],seed[3363],seed[950],seed[943],seed[782],seed[605],seed[1028],seed[2523],seed[183],seed[2348],seed[3392],seed[2437],seed[2244],seed[3496],seed[3128],seed[3248],seed[3970],seed[322],seed[261],seed[180],seed[481],seed[74],seed[4001],seed[2185],seed[1967],seed[1195],seed[1192],seed[2184],seed[1332],seed[788],seed[3270],seed[2533],seed[3762],seed[3870],seed[1563],seed[1226],seed[1276],seed[3533],seed[4020],seed[749],seed[218],seed[4010],seed[3005],seed[2080],seed[862],seed[1399],seed[405],seed[1131],seed[1706],seed[3911],seed[2912],seed[417],seed[3475],seed[3537],seed[369],seed[1765],seed[3010],seed[3967],seed[3028],seed[2595],seed[1802],seed[1172],seed[3075],seed[4059],seed[371],seed[1145],seed[2299],seed[1745],seed[2411],seed[3587],seed[277],seed[2481],seed[479],seed[2574],seed[3662],seed[1531],seed[1323],seed[2720],seed[3286],seed[555],seed[3750],seed[2302],seed[3746],seed[3882],seed[3143],seed[2116],seed[821],seed[2748],seed[2821],seed[1352],seed[1512],seed[1129],seed[1496],seed[43],seed[2710],seed[1891],seed[2225],seed[2841],seed[4014],seed[1998],seed[3801],seed[264],seed[1360],seed[1173],seed[1081],seed[273],seed[1290],seed[3411],seed[399],seed[182],seed[651],seed[3930],seed[2043],seed[314],seed[999],seed[1777],seed[3806],seed[1959],seed[3855],seed[186],seed[3193],seed[857],seed[3251],seed[2275],seed[2854],seed[3182],seed[3996],seed[1047],seed[3839],seed[978],seed[2757],seed[968],seed[1054],seed[1536],seed[3730],seed[3227],seed[1449],seed[3512],seed[2618],seed[2147],seed[3300],seed[2284],seed[1826],seed[2454],seed[305],seed[2916],seed[378],seed[738],seed[2745],seed[2815],seed[3266],seed[2246],seed[1717],seed[1311],seed[3452],seed[1660],seed[3168],seed[3416],seed[2218],seed[3641],seed[3710],seed[3895],seed[1893],seed[3057],seed[1964],seed[2782],seed[3539],seed[1614],seed[94],seed[3199],seed[2006],seed[1196],seed[116],seed[4046],seed[3958],seed[2946],seed[3777],seed[4069],seed[3650],seed[1317],seed[3279],seed[3986],seed[2221],seed[629],seed[485],seed[2562],seed[3337],seed[2696],seed[2151],seed[1072],seed[2753],seed[2001],seed[1672],seed[401],seed[221],seed[764],seed[3447],seed[3657],seed[2473],seed[2769],seed[5],seed[2883],seed[2892],seed[1730],seed[3485],seed[2358],seed[735],seed[3589],seed[1457],seed[3955],seed[2176],seed[3542],seed[197],seed[1204],seed[1969],seed[1374],seed[2292],seed[3984],seed[627],seed[577],seed[3766],seed[316],seed[3681],seed[2903],seed[1477],seed[1393],seed[2138],seed[3090],seed[4051],seed[2182],seed[2103],seed[2694],seed[1709],seed[2444],seed[1671],seed[2127],seed[3885],seed[3486],seed[2713],seed[2251],seed[1798],seed[3360],seed[988],seed[159],seed[926],seed[3034],seed[849],seed[2861],seed[4049],seed[2553],seed[476],seed[2156],seed[573],seed[145],seed[304],seed[3051],seed[956],seed[704],seed[174],seed[1159],seed[1902],seed[3577],seed[1699],seed[920],seed[911],seed[1067],seed[1168],seed[3756],seed[1112],seed[255],seed[622],seed[2441],seed[1681],seed[1342],seed[3894],seed[3856],seed[105],seed[1189],seed[3302],seed[2943],seed[3946],seed[2404],seed[2989],seed[565],seed[699],seed[923],seed[263],seed[1643],seed[3272],seed[2197],seed[1139],seed[2525],seed[3097],seed[1492],seed[3659],seed[1467],seed[670],seed[1823],seed[634],seed[1101],seed[191],seed[1381],seed[3289],seed[2427],seed[3281],seed[3440],seed[3303],seed[1750],seed[2440],seed[2693],seed[1238],seed[3370],seed[2093],seed[884],seed[773],seed[784],seed[3732],seed[78],seed[3778],seed[1202],seed[1971],seed[3961],seed[179],seed[3022],seed[297],seed[2934],seed[2742],seed[1795],seed[684],seed[2935],seed[2457],seed[2798],seed[2049],seed[903],seed[18],seed[3860],seed[1504],seed[1723],seed[2991],seed[1309],seed[2099],seed[3615],seed[3943],seed[1205],seed[3886],seed[3085],seed[2399],seed[2464],seed[2126],seed[797],seed[1090],seed[3245],seed[2121],seed[146],seed[3887],seed[976],seed[115],seed[861],seed[2035],seed[955],seed[1338],seed[614],seed[3497],seed[2367],seed[1843],seed[1888],seed[1876],seed[1575],seed[3335],seed[1383],seed[1208],seed[1216],seed[3350],seed[1108],seed[1503],seed[3724],seed[3872],seed[294],seed[836],seed[706],seed[2010],seed[1160],seed[3479],seed[2304],seed[790],seed[1017],seed[440],seed[4057],seed[2548],seed[474],seed[582],seed[2328],seed[2783],seed[3186],seed[2175],seed[1014],seed[2293],seed[1701],seed[887],seed[3989],seed[2253],seed[2867],seed[1137],seed[2990],seed[3118],seed[3261],seed[1578],seed[2613],seed[1475],seed[649],seed[2590],seed[656],seed[827],seed[1435],seed[1490],seed[1919],seed[353],seed[3201],seed[1863],seed[2177],seed[2965],seed[3393],seed[3742],seed[775],seed[2429],seed[1735],seed[1976],seed[2270],seed[1120],seed[325],seed[592],seed[3365],seed[916],seed[2592],seed[647],seed[2298],seed[3857],seed[2586],seed[894],seed[1494],seed[47],seed[2104],seed[2708],seed[2929],seed[3383],seed[162],seed[1165],seed[2289],seed[3030],seed[433],seed[4025],seed[323],seed[1178],seed[3442],seed[1821],seed[276],seed[4058],seed[1769],seed[740],seed[2305],seed[4030],seed[3660],seed[3796],seed[1083],seed[2608],seed[2852],seed[2770],seed[743],seed[3607],seed[1417],seed[36],seed[202],seed[3202],seed[2220],seed[3269],seed[1087],seed[268],seed[707],seed[1171],seed[2597],seed[92],seed[2800],seed[1235],seed[638],seed[1355],seed[472],seed[772],seed[501],seed[224],seed[1977],seed[3980],seed[1591],seed[946],seed[3709],seed[2313],seed[3928],seed[2276],seed[3080],seed[4043],seed[1647],seed[1240],seed[2067],seed[62],seed[1772],seed[3686],seed[2066],seed[3890],seed[2976],seed[1625],seed[144],seed[2317],seed[2306],seed[3902],seed[3617],seed[1203],seed[3819],seed[3361],seed[135],seed[67],seed[2986],seed[583],seed[79],seed[2310],seed[3956],seed[3752],seed[3760],seed[3025],seed[3287],seed[2308],seed[818],seed[2507],seed[2765],seed[2759],seed[2729],seed[2352],seed[2274],seed[1088],seed[3165],seed[1537],seed[2402],seed[2476],seed[2530],seed[3521],seed[381],seed[2278],seed[3],seed[3152],seed[3763],seed[3206],seed[2637],seed[3222],seed[2674],seed[538],seed[1057],seed[3735],seed[3805],seed[260],seed[2071],seed[3765],seed[567],seed[3802],seed[3768],seed[2107],seed[1678],seed[3726],seed[3111],seed[3784],seed[10],seed[2911],seed[2227],seed[2233],seed[2871],seed[231],seed[1903],seed[3119],seed[1130],seed[2921],seed[3472],seed[2144],seed[3861],seed[3618],seed[1652],seed[3487],seed[2164],seed[2747],seed[1937],seed[2763],seed[2682],seed[3842],seed[598],seed[3716],seed[2996],seed[2020],seed[2417],seed[1636],seed[1307],seed[3653],seed[2688],seed[3776],seed[1605],seed[3788],seed[111],seed[3545],seed[674],seed[3336],seed[3547],seed[3863],seed[1147],seed[451],seed[1291],seed[1434],seed[3780],seed[985],seed[2413],seed[505],seed[522],seed[364],seed[1308],seed[3164],seed[3978],seed[4036],seed[2393],seed[3058],seed[2834],seed[632],seed[3810],seed[3525],seed[1713],seed[2593],seed[913],seed[2450],seed[3783],seed[2646],seed[2802],seed[1901],seed[2610],seed[2259],seed[2432],seed[2790],seed[3723],seed[166],seed[1297],seed[2909],seed[2754],seed[3546],seed[3619],seed[1016],seed[912],seed[1710],seed[981],seed[3439],seed[1414],seed[2543],seed[1190],seed[925],seed[816],seed[243],seed[2055],seed[825],seed[4031],seed[1658],seed[123],seed[3912],seed[686],seed[45],seed[2522],seed[82],seed[219],seed[2860],seed[558],seed[2390],seed[940],seed[217],seed[332],seed[1554],seed[3390],seed[1508],seed[1613],seed[3927],seed[3278],seed[138],seed[2069],seed[1965],seed[3285],seed[963],seed[4005],seed[3434],seed[2849],seed[3817],seed[2621],seed[90],seed[3437],seed[2125],seed[2262],seed[377],seed[2200],seed[3296],seed[2050],seed[4000],seed[132],seed[3596],seed[1657],seed[4093],seed[3744],seed[2307],seed[2953],seed[2162],seed[3637],seed[2247],seed[3157],seed[1814],seed[24],seed[708],seed[2704],seed[1181],seed[2836],seed[1993],seed[3921],seed[59],seed[4055],seed[1033],seed[1128],seed[3065],seed[2799],seed[2158],seed[3459],seed[2409],seed[1320],seed[1945],seed[2650],seed[3652],seed[3638],seed[4012],seed[1753],seed[2607],seed[1683],seed[612],seed[3140],seed[543],seed[3484],seed[1514],seed[524],seed[2531],seed[2668],seed[1861],seed[1187],seed[609],seed[1346],seed[1126],seed[2947],seed[1053],seed[2179],seed[3673],seed[3597],seed[1906],seed[712],seed[1687],seed[3061],seed[530],seed[19],seed[2766],seed[3282],seed[2920],seed[3430],seed[2949],seed[1348],seed[844],seed[1201],seed[838],seed[2029],seed[2466],seed[1925],seed[3888],seed[3339],seed[2436],seed[455],seed[553],seed[1365],seed[1640],seed[1896],seed[1905],seed[1871],seed[3883],seed[2534],seed[2418],seed[3062],seed[1132],seed[3257],seed[1862],seed[3899],seed[3076],seed[2395],seed[52],seed[3462],seed[1102],seed[3158],seed[3571],seed[3683],seed[1283],seed[1689],seed[3183],seed[1227],seed[2647],seed[3833],seed[288],seed[747],seed[2122],seed[2829],seed[2738],seed[1432],seed[3591],seed[2699],seed[3056],seed[2890],seed[3593],seed[2510],seed[2297],seed[1106],seed[2282],seed[2456],seed[477],seed[3297],seed[2728],seed[345],seed[2271],seed[3029],seed[3457],seed[2767],seed[1061],seed[1140],seed[107],seed[3268],seed[3351],seed[289],seed[100],seed[930],seed[678],seed[2888],seed[88],seed[1279],seed[1464],seed[2709],seed[1186],seed[1161],seed[2167],seed[1143],seed[3914],seed[2971],seed[3654],seed[2128],seed[2975],seed[1935],seed[2505],seed[3785],seed[1078],seed[2028],seed[1724],seed[91],seed[3469],seed[1560],seed[3079],seed[2814],seed[2707],seed[315],seed[414],seed[3612],seed[3506],seed[860],seed[1956],seed[3749],seed[1595],seed[1095],seed[1736],seed[786],seed[338],seed[56],seed[2420],seed[902],seed[504],seed[129],seed[3362],seed[1242],seed[3397],seed[1448],seed[2111],seed[3731],seed[2733],seed[4090],seed[2149],seed[3556],seed[3689],seed[1799],seed[2740],seed[1409],seed[2558],seed[1879],seed[1887],seed[2286],seed[3532],seed[2141],seed[1287],seed[3616],seed[1587],seed[939],seed[3705],seed[3694],seed[702],seed[2915],seed[42],seed[1326],seed[3908],seed[1356],seed[223],seed[868],seed[2686],seed[3418],seed[3324],seed[4065],seed[204],seed[2132],seed[2488],seed[2662],seed[2007],seed[2692],seed[1113],seed[1426],seed[3600],seed[3864],seed[12],seed[2596],seed[70],seed[2046],seed[3332],seed[2135],seed[636],seed[980],seed[2098],seed[3918],seed[619],seed[2204],seed[1149],seed[390],seed[1986],seed[3410],seed[1405],seed[2567],seed[1616],seed[2508],seed[3117],seed[3661],seed[1727],seed[1661],seed[3059],seed[3255],seed[533],seed[2323],seed[502],seed[2446],seed[3129],seed[842],seed[1872],seed[2169],seed[1921],seed[1382],seed[2619],seed[2287],seed[1366],seed[2906],seed[3413],seed[576],seed[3929],seed[1979],seed[1465],seed[3502],seed[1809],seed[3432],seed[3323],seed[2605],seed[2573],seed[357],seed[630],seed[3798],seed[3540],seed[427],seed[2572],seed[1371],seed[669],seed[2524],seed[3233],seed[1251],seed[2261],seed[407],seed[3877],seed[4013],seed[723],seed[2166],seed[854],seed[635],seed[3223],seed[3687],seed[2474],seed[256],seed[1237],seed[1629],seed[1631],seed[834],seed[3012],seed[1786],seed[1819],seed[2335],seed[1856],seed[3315],seed[134],seed[1328],seed[2559],seed[3625],seed[4039],seed[886],seed[713],seed[1731],seed[2615],seed[1599],seed[1091],seed[318],seed[3960],seed[410],seed[2114],seed[1122],seed[2130],seed[3874],seed[1573],seed[863],seed[3124],seed[2571],seed[2239],seed[450],seed[785],seed[4],seed[3713],seed[3519],seed[965],seed[3628],seed[239],seed[2865],seed[1150],seed[3633],seed[673],seed[2891],seed[2431],seed[2015],seed[120],seed[2374],seed[1991],seed[2497],seed[663],seed[2058],seed[1547],seed[334],seed[3103],seed[233],seed[2653],seed[2490],seed[828],seed[648],seed[896],seed[3349],seed[1583],seed[789],seed[3375],seed[3120],seed[3342],seed[534],seed[3741],seed[3682],seed[383],seed[2514],seed[3037],seed[645],seed[3108],seed[3247],seed[2962],seed[1598],seed[2599],seed[3088],seed[3169],seed[1927],seed[3624],seed[1722],seed[208],seed[1422],seed[1153],seed[3027],seed[2148],seed[1728],seed[1637],seed[3516],seed[1110],seed[1559],seed[3923],seed[2846],seed[588],seed[4092],seed[570],seed[2521],seed[3275],seed[2520],seed[199],seed[2551],seed[2192],seed[1146],seed[556],seed[1674],seed[744],seed[2294],seed[3074],seed[1104],seed[2835],seed[1258],seed[388],seed[979],seed[545],seed[1663],seed[2252],seed[2318],seed[719],seed[2874],seed[4073],seed[2687],seed[3853],seed[3004],seed[3319],seed[2830],seed[280],seed[1200],seed[2651],seed[1176],seed[38],seed[185],seed[3376],seed[3477],seed[1483],seed[2248],seed[2109],seed[1865],seed[858],seed[4045],seed[3811],seed[3053],seed[1357],seed[660],seed[3288],seed[2459],seed[3603],seed[2034],seed[1164],seed[2760],seed[2701],seed[1797],seed[914],seed[3252],seed[4076],seed[2052],seed[235],seed[2316],seed[3972],seed[1949],seed[3913],seed[2054],seed[1783],seed[599],seed[3399],seed[3114],seed[99],seed[1314],seed[847],seed[2914],seed[3561],seed[3708],seed[1516],seed[490],seed[2718],seed[17],seed[595],seed[701],seed[26],seed[1923],seed[2414],seed[1368],seed[2353],seed[3953],seed[1827],seed[2272],seed[3283],seed[3954],seed[757],seed[953],seed[561],seed[178],seed[1733],seed[3535],seed[2356],seed[3292],seed[61],seed[574],seed[1519],seed[2372],seed[3271],seed[590],seed[1794],seed[2664],seed[1756],seed[3718],seed[3344],seed[1911],seed[1789],seed[1751],seed[1719],seed[3728],seed[3588],seed[1900],seed[2797],seed[724],seed[1438],seed[4075],seed[475],seed[3425],seed[1300],seed[681],seed[813],seed[3256],seed[2207],seed[1757],seed[2758],seed[3017],seed[3389],seed[3523],seed[1339],seed[3396],seed[520],seed[136],seed[1768],seed[3348],seed[3733],seed[3013],seed[3384],seed[1858],seed[1424],seed[2764],seed[2375],seed[2925],seed[2931],seed[1655],seed[1466],seed[3629],seed[2076],seed[1749],seed[148],seed[3951],seed[1032],seed[426],seed[2471],seed[34],seed[2667],seed[3039],seed[2630],seed[537],seed[2101],seed[1386],seed[2256],seed[594],seed[4053],seed[3636],seed[375],seed[1479],seed[1632],seed[1505],seed[3826],seed[1961],seed[1646],seed[2863],seed[1299],seed[229],seed[3455],seed[855],seed[2509],seed[780],seed[616],seed[1779],seed[3721],seed[2695],seed[1040],seed[1407],seed[3920],seed[626],seed[319],seed[871],seed[164],seed[2008],seed[3042],seed[1058],seed[3020],seed[2979],seed[3041],seed[3906],seed[1350],seed[984],seed[2542],seed[3809],seed[951],seed[2243],seed[889],seed[1079],seed[734],seed[3670],seed[2478],seed[3676],seed[3568],seed[3184],seed[3595],seed[3083],seed[434],seed[275],seed[1851],seed[4009],seed[819],seed[736],seed[3758],seed[3774],seed[1952],seed[1897],seed[2153],seed[1633],seed[2545],seed[3761],seed[3449],seed[907],seed[1524],seed[2194],seed[2967],seed[549],seed[2649],seed[1343],seed[2344],seed[1228],seed[2685],seed[1972],seed[1545],seed[2266],seed[3294],seed[2658],seed[809],seed[2094],seed[2363],seed[1796],seed[3702],seed[2455],seed[1468],seed[3189],seed[1572],seed[2584],seed[2462],seed[142],seed[812],seed[1517],seed[2812],seed[814],seed[1840],seed[1018],seed[2461],seed[3696],seed[3706],seed[1580],seed[503],seed[1764],seed[802],seed[1626],seed[1315],seed[2143],seed[3379],seed[2952],seed[2406],seed[2671],seed[3318],seed[3747],seed[2235],seed[3828],seed[3264],seed[1369],seed[3854],seed[1493],seed[3720],seed[3808],seed[1020],seed[3087],seed[1260],seed[3021],seed[3795],seed[1319],seed[328],seed[2351],seed[877],seed[1568],seed[3018],seed[1335],seed[1985],seed[1557],seed[2722],seed[193],seed[498],seed[3427],seed[2228],seed[600],seed[2850],seed[3064],seed[1778],seed[207],seed[363],seed[449],seed[3215],seed[4048],seed[1246],seed[1914],seed[4027],seed[3896],seed[4023],seed[413],seed[2036],seed[562],seed[1313],seed[2743],seed[2097],seed[1695],seed[141],seed[3668],seed[966],seed[33],seed[1141],seed[2350],seed[1834],seed[3259],seed[737],seed[2828],seed[547],seed[1274],seed[2768],seed[2453],seed[3214],seed[2477],seed[883],seed[3719],seed[2908],seed[1780],seed[1673],seed[29],seed[2540],seed[3693],seed[3498],seed[1004],seed[3737],seed[2755],seed[2676],seed[1446],seed[484],seed[1922],seed[3038],seed[339],seed[792],seed[2697],seed[4091],seed[2794],seed[3408],seed[3395],seed[535],seed[3775],seed[3078],seed[1878],seed[3356],seed[1530],seed[2236],seed[3309],seed[526],seed[841],seed[2725],seed[650],seed[3197],seed[3821],seed[2472],seed[2095],seed[687],seed[1670],seed[2726],seed[658],seed[948],seed[575],seed[3916],seed[2493],seed[2938],seed[2030],seed[2875],seed[4029],seed[3422],seed[3889],seed[3273],seed[1742],seed[3131],seed[222],seed[2019],seed[3474],seed[3634],seed[2386],seed[1125],seed[3651],seed[3156],seed[927],seed[606],seed[2555],seed[941],seed[2869],seed[3398],seed[1828],seed[1607],seed[2864],seed[1296],seed[905],seed[1940],seed[2154],seed[3196],seed[2354],seed[3979],seed[303],seed[3443],seed[1292],seed[1423],seed[4034],seed[3580],seed[3552],seed[2910],seed[2403],seed[4032],seed[1784],seed[1071],seed[327],seed[3132],seed[3663],seed[2012],seed[1413],seed[3448],seed[1182],seed[3941],seed[3191],seed[3602],seed[3254],seed[329],seed[2378],seed[2070],seed[1213],seed[3126],seed[1712],seed[3170],seed[3220],seed[717],seed[910],seed[2504],seed[1249],seed[3490],seed[691],seed[3262],seed[3656],seed[1523],seed[237],seed[1609],seed[837],seed[1581],seed[1838],seed[1043],seed[2749],seed[1877],seed[3782],seed[1837],seed[1930],seed[1694],seed[3428],seed[2330],seed[3583],seed[1388],seed[487],seed[1170],seed[2626],seed[869],seed[2326],seed[2032],seed[1848],seed[2479],seed[171],seed[2113],seed[1391],seed[348],seed[2882],seed[1617],seed[3697],seed[175],seed[1770],seed[3831],seed[897],seed[2907],seed[28],seed[1135],seed[3423],seed[102],seed[731],seed[2784],seed[2380],seed[2970],seed[2904],seed[1015],seed[3692],seed[1918],seed[2617],seed[2206],seed[402],seed[2632],seed[1100],seed[803],seed[165],seed[1886],seed[2727],seed[853],seed[3293],seed[685],seed[2347],seed[3844],seed[2215],seed[1076],seed[124],seed[1118],seed[720],seed[415],seed[508],seed[1615],seed[3301],seed[1261],seed[4007],seed[3959],seed[3703],seed[2640],seed[2536],seed[2622],seed[895],seed[1544],seed[40],seed[1232],seed[1373],seed[2312],seed[98],seed[935],seed[254],seed[1853],seed[1939],seed[2778],seed[3135],seed[3530],seed[832],seed[721],seed[3380],seed[2336],seed[431],seed[3372],seed[77],seed[2415],seed[1608],seed[3401],seed[3868],seed[480],seed[1041],seed[1295],seed[3331],seed[152],seed[711],seed[1639],seed[72],seed[960],seed[2387],seed[3509],seed[845],seed[3992],seed[2995],seed[970],seed[3926],seed[3225],seed[1395],seed[3415],seed[2423],seed[4033],seed[2937],seed[901],seed[1589],seed[3195],seed[1324],seed[3977],seed[2240],seed[3579],seed[1577],seed[1996],seed[3609],seed[1570],seed[1535],seed[2872],seed[3901],seed[810],seed[4060],seed[75],seed[932],seed[3329],seed[625],seed[856],seed[2222],seed[2343],seed[2059],seed[3759],seed[1430],seed[2974],seed[460],seed[2405],seed[2661],seed[4002],seed[1664],seed[2408],seed[416],seed[1055],seed[1436],seed[389],seed[3304],seed[3123],seed[2998],seed[1501],seed[3263],seed[4087],seed[3938],seed[2443],seed[2340],seed[1298],seed[1542],seed[794],seed[380],seed[1488],seed[1656],seed[548],seed[1451],seed[1973],seed[2893],seed[640],seed[3134],seed[3932],seed[3613],seed[2416],seed[3518],seed[1217],seed[3127],seed[343],seed[540],seed[2837],seed[2048],seed[257],seed[3404],seed[302],seed[65],seed[804],seed[1119],seed[2484],seed[3818],seed[2988],seed[2022],seed[1481],seed[489],seed[3374],seed[2897],seed[1364],seed[2021],seed[2535],seed[992],seed[1269],seed[2956],seed[993],seed[1460],seed[1994],seed[3646],seed[3834],seed[1321],seed[441],seed[1404],seed[2039],seed[791],seed[103],seed[3113],seed[3995],seed[362],seed[2072],seed[3631],seed[311],seed[3517],seed[2460],seed[3274],seed[1932],seed[2657],seed[891],seed[446],seed[1392],seed[3205],seed[3966],seed[1500],seed[3569],seed[3876],seed[2499],seed[1708],seed[1836],seed[1690],seed[2933],seed[32],seed[2680],seed[866],seed[1686],seed[2684],seed[513],seed[2161],seed[3866],seed[2614],seed[1134],seed[3063],seed[517],seed[921],seed[3298],seed[1995],seed[2005],seed[1476],seed[3325],seed[2842],seed[3804],seed[3414],seed[3204],seed[97],seed[1486],seed[922],seed[3240],seed[1233],seed[117],seed[1803],seed[807],seed[3492],seed[3310],seed[709],seed[2320],seed[1484],seed[2873],seed[1805],seed[2321],seed[2364],seed[1954],seed[1926],seed[1532],seed[4095],seed[2537],seed[3016],seed[727],seed[1459],seed[1241],seed[2868],seed[4068],seed[2856],seed[1285],seed[430],seed[1635],seed[2018],seed[621],seed[2969],seed[2234],seed[661],seed[2376],seed[1820],seed[945],seed[3865],seed[2425],seed[1303],seed[1624],seed[2331],seed[3420],seed[2024],seed[2000],seed[739],seed[1791],seed[3322],seed[1641],seed[283],seed[3534],seed[3549],seed[1738],seed[1390],seed[1062],seed[1450],seed[1539],seed[187],seed[2337],seed[1763],seed[1385],seed[406],seed[958],seed[2663],seed[688],seed[551],seed[2160],seed[2397],seed[589],seed[372],seed[1021],seed[1978],seed[689],seed[39],seed[2918],seed[55],seed[1497],seed[3513],seed[2612],seed[11],seed[2641],seed[677],seed[1329],seed[3983],seed[3666],seed[1097],seed[21],seed[3942],seed[1225],seed[301],seed[1243],seed[3105],seed[2419],seed[1431],seed[2196],seed[3444],seed[1666],seed[1868],seed[2051],seed[1133],seed[463],seed[3489],seed[808],seed[1928],seed[4088],seed[1529],seed[3308],seed[292],seed[2756],seed[425],seed[2655],seed[698],seed[1439],seed[633],seed[3655],seed[1412],seed[1920],seed[2487],seed[149],seed[2213],seed[93],seed[1885],seed[211],seed[2085],seed[3559],seed[3066],seed[1157],seed[2624],seed[266],seed[2566],seed[1792],seed[1755],seed[982],seed[4089],seed[7],seed[2642],seed[1693],seed[1725],seed[2838],seed[1001],seed[1654],seed[2065],seed[3473],seed[3213],seed[1705],seed[2702],seed[1194],seed[783],seed[1094],seed[2277],seed[1951],seed[157],seed[885],seed[1600],seed[3216],seed[3321],seed[1844],seed[3077],seed[2332],seed[3647],seed[2057],seed[1565],seed[833],seed[3386],seed[3779],seed[3433],seed[3903],seed[2635],seed[1815],seed[2594],seed[2656],seed[665],seed[541],seed[3727],seed[3584],seed[3755],seed[3508],seed[4079],seed[3878],seed[3981],seed[615],seed[664],seed[766],seed[1254],seed[3642],seed[271],seed[2470],seed[3226],seed[3159],seed[1869],seed[1188],seed[779],seed[733],seed[2383],seed[942],seed[2482],seed[3851],seed[3799],seed[801],seed[3910],seed[2163],seed[3846],seed[618],seed[467],seed[3424],seed[3892],seed[2698],seed[1831],seed[512],seed[2880],seed[3050],seed[1267],seed[585],seed[3820],seed[3234],seed[3852],seed[3740],seed[3585],seed[872],seed[1331],seed[203],seed[557],seed[6],seed[1966],seed[3950],seed[2993],seed[3160],seed[2042],seed[1376],seed[31],seed[110],seed[1253],seed[3684],seed[195],seed[1069],seed[820],seed[287],seed[795],seed[1622],seed[13],seed[421],seed[3369],seed[3291],seed[2279],seed[671],seed[3897],seed[971],seed[3095],seed[987],seed[2819],seed[4037],seed[3092],seed[1312],seed[1334],seed[2463],seed[3040],seed[1944],seed[3531],seed[1669],seed[3503],seed[1592],seed[2014],seed[3594],seed[458],seed[3526],seed[776],seed[1304],seed[1857],seed[365],seed[2371],seed[2538],seed[1787],seed[478],seed[3945],seed[1515],seed[358],seed[796],seed[2980],seed[2775],seed[1782],seed[2576],seed[1219],seed[3840],seed[459],seed[3949],seed[3099],seed[3149],seed[3347],seed[1419],seed[2291],seed[2807],seed[2583],seed[3807],seed[2737],seed[4086],seed[683],seed[563],seed[1220],seed[3622],seed[2091],seed[2361],seed[1845],seed[2515],seed[4042],seed[2940],seed[176],seed[514],seed[2031],seed[2627],seed[1586],seed[2564],seed[4015],seed[3773],seed[623],seed[1566],seed[1543],seed[423],seed[497],seed[3674],seed[2117],seed[2193],seed[1754],seed[2879],seed[2480],seed[560],seed[1638],seed[1082],seed[3501],seed[3054],seed[300],seed[1847],seed[3144],seed[2691],seed[3212],seed[2550],seed[2195],seed[1527],seed[781],seed[3453],seed[4016],seed[121],seed[2392],seed[793],seed[753],seed[1433],seed[2496],seed[1175],seed[2285],seed[591],seed[1711],seed[3743],seed[212],seed[1103],seed[360],seed[3825],seed[4061],seed[2498],seed[1953],seed[750],seed[2957],seed[2889],seed[1256],seed[3769],seed[3880],seed[3848],seed[216],seed[1471],seed[1620],seed[3898],seed[2845],seed[2881],seed[3190],seed[1347],seed[1401],seed[1833],seed[3841],seed[2774],seed[4019],seed[1415],seed[694],seed[2506],seed[1049],seed[3174],seed[2930],seed[1759],seed[2366],seed[3794],seed[1470],seed[214],seed[404],seed[777],seed[3873],seed[1367],seed[3973],seed[3468],seed[242],seed[3265],seed[1507],seed[654],seed[3177],seed[409],seed[1025],seed[22],seed[986],seed[607],seed[1406],seed[3176],seed[2438],seed[2365],seed[104],seed[2791],seed[2750],seed[2083],seed[48],seed[225],seed[1692],seed[787],seed[2955],seed[1281],seed[3280],seed[3757],seed[3081],seed[3627],seed[3738],seed[3239],seed[1904],seed[2926],seed[3210],seed[3388],seed[3172],seed[1700],seed[2703],seed[2037],seed[1474],seed[1734],seed[1289],seed[1518],seed[2381],seed[1999],seed[1988],seed[1950],seed[2611],seed[597],seed[3464],seed[3748],seed[96],seed[3217],seed[1068],seed[1003],seed[1597],seed[973],seed[3522],seed[246],seed[878],seed[278],seed[904],seed[2789],seed[2665],seed[3002],seed[3753],seed[370],seed[2136],seed[393],seed[2424],seed[1525],seed[2556],seed[438],seed[1379],seed[113],seed[1548],seed[934],seed[3704],seed[2502],seed[1648],seed[1808],seed[1051],seed[2301],seed[758],seed[2217],seed[3793],seed[1807],seed[3070],seed[937],seed[2721],seed[2013],seed[2866],seed[725],seed[3491],seed[3644],seed[1506],seed[1013],seed[4035],seed[3871],seed[1612],seed[2963],seed[240],seed[20],seed[1601],seed[3564],seed[3402],seed[933],seed[3900],seed[1567],seed[1098],seed[1721],seed[2648],seed[385],seed[2486],seed[3480],seed[774],seed[3739],seed[2339],seed[3515],seed[1322],seed[3218],seed[2853],seed[2932],seed[2255],seed[2673],seed[752],seed[188],seed[1375],seed[58],seed[1060],seed[3368],seed[73],seed[147],seed[3707],seed[639],seed[1582],seed[326],seed[4081],seed[230],seed[2981],seed[2512],seed[445],seed[471],seed[4066],seed[2483],seed[2820],seed[3639],seed[299],seed[3466],seed[3091],seed[2563],seed[2539],seed[1163],seed[715],seed[308],seed[184],seed[2554],seed[569],seed[2400],seed[2825],seed[1907],seed[1746],seed[2549],seed[64],seed[51],seed[1027],seed[2785],seed[3745],seed[566],seed[2439],seed[190],seed[1183],seed[2643],seed[4028],seed[601],seed[466],seed[995],seed[3791],seed[2964],seed[2090],seed[3700],seed[2303],seed[2449],seed[2818],seed[2033],seed[68],seed[2788],seed[2810],seed[2341],seed[2263],seed[1358],seed[2142],seed[2283],seed[2370],seed[1007],seed[1943],seed[464],seed[3451],seed[716],seed[3044],seed[1982],seed[352],seed[2190],seed[2919],seed[2858],seed[2045],seed[295],seed[2202],seed[2811],seed[3614],seed[2448],seed[3813],seed[2009],seed[3026],seed[2334],seed[1980],seed[432],seed[1957],seed[2848],seed[703],seed[3277],seed[3417],seed[2809],seed[3109],seed[335],seed[578],seed[2839],seed[1234],seed[1958],seed[3688],seed[1619],seed[1491],seed[3714],seed[652],seed[2081],seed[2659],seed[1302],seed[2532],seed[1114],seed[3884],seed[3907],seed[3536],seed[3258],seed[2369],seed[1551],seed[2744],seed[961],seed[1775],seed[1093],seed[1810],seed[2112],seed[3244],seed[2500],seed[439],seed[653],seed[962],seed[4094],seed[1282],seed[1398],seed[3554],seed[3771],seed[1801],seed[1073],seed[1850],seed[2152],seed[3905],seed[2859],seed[852],seed[2951],seed[3789],seed[1852],seed[1354],seed[1402],seed[3985],seed[2394],seed[1817],seed[2115],seed[1790],seed[3729],seed[2106],seed[2422],seed[1036],seed[150],seed[2973],seed[2273],seed[2064],seed[521],seed[2706],seed[919],seed[641],seed[2016],seed[3881],seed[2541],seed[2519],seed[192],seed[3699],seed[1229],seed[1045],seed[2844],seed[2079],seed[130],seed[546],seed[44],seed[1691],seed[2945],seed[2100],seed[3148],seed[1151],seed[3326],seed[3232],seed[4054],seed[1830],seed[2779],seed[2389],seed[2773],seed[3161],seed[830],seed[2155],seed[2634],seed[696],seed[2966],seed[1121],seed[321],seed[515],seed[550],seed[3314],seed[3320],seed[2178],seed[1248],seed[879],seed[1169],seed[2384],seed[1716],seed[732],seed[3832],seed[1955],seed[1942],seed[949],seed[3922],seed[1881],seed[1854],seed[3429],seed[2205],seed[2445],seed[668],seed[584],seed[1340],seed[1469],seed[646],seed[2],seed[1265],seed[586],seed[3024],seed[2345],seed[2513],seed[8],seed[437],seed[2762],seed[882],seed[1380],seed[108],seed[2265],seed[3999],seed[1806],seed[2752],seed[1191],seed[1009],seed[1344],seed[751],seed[3470],seed[679],seed[2435],seed[398],seed[3231],seed[3338],seed[2985],seed[1992],seed[867],seed[2652],seed[1447],seed[3601],seed[400],seed[2771],seed[2296],seed[2817],seed[3611],seed[2229],seed[3514],seed[3052],seed[1038],seed[210],seed[1325],seed[3988],seed[2060],seed[3667],seed[2560],seed[1704],seed[3575],seed[457],seed[1223],seed[2250],seed[109],seed[3691],seed[1534],seed[2264],seed[523],seed[1099],seed[140],seed[2077],seed[54],seed[2187],seed[3290],seed[697],seed[1762],seed[3645],seed[392],seed[865],seed[2994],seed[1875],seed[241],seed[1330],seed[291],seed[3203],seed[3800],seed[906],seed[3630],seed[2047],seed[14],seed[888],seed[3909],seed[3327],seed[544],seed[3476],seed[3316],seed[1618],seed[1747],seed[2150],seed[158],seed[1277],seed[2732],seed[3071],seed[1372],seed[2672],seed[3493],seed[1662],seed[2430],seed[532],seed[247],seed[1924],seed[3299],seed[2407],seed[1389],seed[2186],seed[2377],seed[1603],seed[3100],seed[3243],seed[3751],seed[1039],seed[4022],seed[3520],seed[2338],seed[1425],seed[331],seed[745],seed[2129],seed[1528],seed[998],seed[3836],seed[3048],seed[447],seed[3426],seed[2442],seed[3971],seed[1306],seed[1034],seed[1895],seed[997],seed[1361],seed[915],seed[2191],seed[3238],seed[422],seed[374],seed[2600],seed[1074],seed[811],seed[2978],seed[373],seed[3764],seed[3933],seed[2644],seed[3675],seed[3610],seed[3671],seed[488],seed[1050],seed[342],seed[3378],seed[2238],seed[2580],seed[2677],seed[817],seed[3359],seed[3006],seed[3093],seed[1744],seed[350],seed[765],seed[3505],seed[2501],seed[1933],seed[3219],seed[611],seed[57],seed[3060],seed[2211],seed[1948],seed[1084],seed[3276],seed[420],seed[469],seed[893],seed[3620],seed[1684],seed[1541],seed[169],seed[1698],seed[1818],seed[1262],seed[2780],seed[344],seed[2902],seed[2581],seed[2620],seed[84],seed[3511],seed[1224],seed[2492],seed[3529],seed[1538],seed[3843],seed[3249],seed[3435],seed[840],seed[2717],seed[3151],seed[2139],seed[351],seed[3236],seed[1884],seed[83],seed[1679],seed[2751],seed[3098],seed[3137],seed[2675],seed[2578],seed[2603],seed[4041],seed[2714],seed[1162],seed[2636],seed[1284],seed[395],seed[419],seed[1177],seed[3106],seed[2958],seed[2568],seed[1011],seed[1048],seed[3551],seed[2203],seed[2491],seed[2922],seed[3538],seed[1136],seed[1070],seed[1677],seed[1456],seed[2041],seed[1630],seed[1198],seed[3094],seed[1623],seed[1936],seed[483],seed[2075],seed[924],seed[1604],seed[3373],seed[1511],seed[2623],seed[468],seed[122],seed[1336],seed[1849],seed[4017],seed[3635],seed[456],seed[3939],seed[657],seed[3450],seed[754],seed[1894],seed[2547],seed[2792],seed[1513],seed[931],seed[1212],seed[2716],seed[2140],seed[3334],seed[3311],seed[3142],seed[2941],seed[1408],seed[3115],seed[1359],seed[672],seed[4006],seed[969],seed[279],seed[2131],seed[368],seed[1030],seed[156],seed[1628],seed[1092],seed[718],seed[3781],seed[2712],seed[2198],seed[1975],seed[262],seed[1584],seed[1761],seed[768],seed[806],seed[1892],seed[1174],seed[296],seed[1855],seed[823],seed[2927],seed[3974],seed[3436],seed[1416],seed[3993],seed[608],seed[2495],seed[3560],seed[2061],seed[3145],seed[1703],seed[2582],seed[3626],seed[1109],seed[1825],seed[2666],seed[511],seed[2281],seed[1318],seed[3850],seed[580],seed[3494],seed[3975],seed[762],seed[2887],seed[2379],seed[349],seed[106],seed[2489],seed[1521],seed[495],seed[1345],seed[3407],seed[2074],seed[778],seed[4084],seed[1167],seed[4021],seed[25],seed[1929],seed[3606],seed[3267],seed[1842],seed[564],seed[2678],seed[1564],seed[2086],seed[1870],seed[2796],seed[3364],seed[403],seed[151],seed[1726],seed[1767],seed[3394],seed[507],seed[2960],seed[1685],seed[3573],seed[1096],seed[572],seed[2451],seed[1288],seed[2209],seed[3623],seed[1962],seed[3672],seed[3228],seed[3400],seed[1832],seed[71],seed[1984],seed[324],seed[376],seed[1555],seed[3211],seed[1916],seed[1378],seed[1215],seed[234],seed[835],seed[881],seed[1042],seed[4024],seed[3237],seed[367],seed[189],seed[3163],seed[2565],seed[1502],seed[3461],seed[967],seed[137],seed[848],seed[1310],seed[2896],seed[282],seed[1873],seed[3454],seed[1989],seed[675],seed[1029],seed[571],seed[496],seed[2087],seed[482],seed[1883],seed[3717],seed[3963],seed[1142],seed[1293],seed[3528],seed[2598],seed[118],seed[1123],seed[3934],seed[742],seed[3504],seed[3133],seed[1561],seed[770],seed[1155],seed[880],seed[2311],seed[2357],seed[1931],seed[4026],seed[3527],seed[1454],seed[700],seed[1180],seed[2426],seed[2781],seed[3406],seed[3815],seed[2241],seed[1341],seed[3162],seed[1675],seed[248],seed[1444],seed[2245],seed[173],seed[170],seed[3701],seed[1247],seed[3665]}),
        .cross_prob(cross_prob),
        .codeword(codeword6),
        .received(received6)
        );
    
    bsc bsc7(
        .clk(clk),
        .reset(reset),
        .seed({seed[426],seed[966],seed[208],seed[2963],seed[2634],seed[283],seed[4017],seed[1315],seed[2560],seed[2387],seed[1724],seed[2509],seed[927],seed[2575],seed[424],seed[2017],seed[1569],seed[3710],seed[1169],seed[2591],seed[2481],seed[1404],seed[874],seed[1491],seed[3883],seed[3967],seed[1599],seed[679],seed[676],seed[1063],seed[2138],seed[2864],seed[2825],seed[2763],seed[3460],seed[2818],seed[1791],seed[13],seed[1196],seed[1111],seed[568],seed[2292],seed[3994],seed[3351],seed[3343],seed[3073],seed[2320],seed[3765],seed[524],seed[3299],seed[3920],seed[2194],seed[1575],seed[3794],seed[1845],seed[2746],seed[3464],seed[3956],seed[3891],seed[1197],seed[2659],seed[2188],seed[1737],seed[2052],seed[1090],seed[1149],seed[2689],seed[652],seed[3328],seed[664],seed[900],seed[3595],seed[1366],seed[3761],seed[3402],seed[429],seed[2175],seed[2394],seed[445],seed[971],seed[1820],seed[736],seed[1098],seed[267],seed[1920],seed[2047],seed[3066],seed[1867],seed[3138],seed[2807],seed[1013],seed[626],seed[476],seed[2432],seed[249],seed[2754],seed[266],seed[3750],seed[151],seed[10],seed[2350],seed[852],seed[3265],seed[388],seed[1973],seed[3881],seed[2772],seed[1461],seed[2023],seed[3076],seed[3263],seed[2495],seed[841],seed[4012],seed[731],seed[138],seed[1236],seed[2987],seed[2336],seed[115],seed[3720],seed[1592],seed[4055],seed[491],seed[313],seed[1322],seed[125],seed[1529],seed[1837],seed[1226],seed[2006],seed[896],seed[2204],seed[372],seed[2829],seed[1494],seed[1789],seed[1877],seed[32],seed[1344],seed[1262],seed[1911],seed[674],seed[3626],seed[435],seed[2528],seed[2161],seed[97],seed[1495],seed[2660],seed[2348],seed[1849],seed[605],seed[3900],seed[3354],seed[3875],seed[997],seed[1385],seed[2847],seed[958],seed[1759],seed[3215],seed[2039],seed[3080],seed[2265],seed[2544],seed[906],seed[3929],seed[908],seed[62],seed[3614],seed[215],seed[2290],seed[4090],seed[2703],seed[3711],seed[3256],seed[164],seed[2679],seed[3851],seed[784],seed[411],seed[2323],seed[507],seed[1654],seed[3936],seed[3529],seed[3544],seed[3637],seed[490],seed[30],seed[2525],seed[837],seed[2124],seed[3541],seed[3699],seed[806],seed[485],seed[1132],seed[3515],seed[1878],seed[1829],seed[4025],seed[329],seed[193],seed[47],seed[203],seed[833],seed[1183],seed[348],seed[3973],seed[2142],seed[3644],seed[2295],seed[1122],seed[2782],seed[3556],seed[2379],seed[452],seed[1295],seed[1524],seed[1434],seed[2501],seed[1472],seed[1025],seed[3426],seed[600],seed[2063],seed[3240],seed[1508],seed[101],seed[1754],seed[2428],seed[2210],seed[1287],seed[3560],seed[1847],seed[1413],seed[393],seed[2885],seed[750],seed[2189],seed[3921],seed[2106],seed[1931],seed[3923],seed[2723],seed[3659],seed[3741],seed[3376],seed[3201],seed[46],seed[3686],seed[179],seed[1022],seed[1717],seed[111],seed[1251],seed[1283],seed[3648],seed[1039],seed[3363],seed[4045],seed[1813],seed[3123],seed[120],seed[683],seed[950],seed[2135],seed[2258],seed[2768],seed[3456],seed[1065],seed[812],seed[3119],seed[486],seed[1840],seed[1305],seed[2624],seed[3554],seed[1555],seed[1081],seed[3919],seed[3386],seed[102],seed[2317],seed[1735],seed[946],seed[2195],seed[409],seed[1456],seed[1546],seed[2452],seed[3745],seed[2122],seed[3910],seed[2959],seed[1469],seed[4086],seed[77],seed[2683],seed[930],seed[3840],seed[471],seed[3014],seed[2526],seed[22],seed[3521],seed[543],seed[3346],seed[3389],seed[1856],seed[1425],seed[1630],seed[140],seed[1726],seed[2310],seed[15],seed[2633],seed[3278],seed[630],seed[2981],seed[1255],seed[3597],seed[487],seed[3121],seed[2519],seed[2248],seed[1821],seed[980],seed[1916],seed[2127],seed[1927],seed[880],seed[168],seed[1693],seed[3410],seed[1384],seed[1954],seed[2021],seed[3028],seed[295],seed[2173],seed[1695],seed[1487],seed[494],seed[3372],seed[2845],seed[1997],seed[1447],seed[2190],seed[621],seed[3530],seed[1083],seed[1522],seed[1317],seed[924],seed[1518],seed[1310],seed[3142],seed[1679],seed[2249],seed[1898],seed[2802],seed[994],seed[234],seed[2433],seed[2618],seed[2539],seed[3668],seed[480],seed[3161],seed[1184],seed[3196],seed[1962],seed[3200],seed[1077],seed[3718],seed[2655],seed[3519],seed[73],seed[823],seed[2030],seed[3436],seed[3226],seed[536],seed[2028],seed[1311],seed[3636],seed[2706],seed[3949],seed[1551],seed[2270],seed[1961],seed[1335],seed[2380],seed[3183],seed[3455],seed[1258],seed[3144],seed[3168],seed[538],seed[3630],seed[3939],seed[3139],seed[3812],seed[1643],seed[2642],seed[2684],seed[1797],seed[3645],seed[2974],seed[1527],seed[3433],seed[3622],seed[651],seed[3173],seed[3228],seed[1026],seed[3442],seed[2403],seed[1362],seed[697],seed[3513],seed[2695],seed[2606],seed[2532],seed[1772],seed[3380],seed[1430],seed[12],seed[1966],seed[391],seed[3242],seed[3109],seed[2546],seed[1218],seed[1652],seed[2923],seed[1059],seed[1783],seed[37],seed[855],seed[527],seed[2902],seed[3866],seed[1155],seed[2469],seed[2031],seed[3983],seed[3149],seed[1386],seed[55],seed[2739],seed[1429],seed[2445],seed[3182],seed[1681],seed[2038],seed[1608],seed[2326],seed[1268],seed[3740],seed[2529],seed[1440],seed[776],seed[2637],seed[1248],seed[1725],seed[444],seed[3486],seed[159],seed[2698],seed[3928],seed[99],seed[1102],seed[1347],seed[3469],seed[3682],seed[1156],seed[1137],seed[1649],seed[3806],seed[1906],seed[4040],seed[2792],seed[2785],seed[1894],seed[2652],seed[3036],seed[3448],seed[3214],seed[3322],seed[2410],seed[814],seed[3338],seed[572],seed[3514],seed[71],seed[2113],seed[2430],seed[3435],seed[2828],seed[3533],seed[3255],seed[2111],seed[1776],seed[1399],seed[2202],seed[1841],seed[1061],seed[2280],seed[2774],seed[1596],seed[3086],seed[2992],seed[2570],seed[2827],seed[3826],seed[1383],seed[3972],seed[3814],seed[1237],seed[525],seed[3795],seed[1094],seed[3859],seed[314],seed[3192],seed[395],seed[530],seed[1744],seed[457],seed[364],seed[2055],seed[3285],seed[3395],seed[1235],seed[1660],seed[1123],seed[1722],seed[518],seed[3027],seed[170],seed[3450],seed[3083],seed[3445],seed[2125],seed[539],seed[341],seed[1870],seed[3500],seed[3403],seed[1680],seed[3416],seed[685],seed[3393],seed[1353],seed[1133],seed[1541],seed[2443],seed[3154],seed[1192],seed[2256],seed[3269],seed[2910],seed[2567],seed[427],seed[540],seed[1532],seed[2158],seed[2631],seed[890],seed[2592],seed[3661],seed[109],seed[942],seed[1479],seed[3052],seed[2473],seed[3522],seed[2468],seed[4093],seed[1459],seed[2770],seed[2565],seed[469],seed[4041],seed[2645],seed[260],seed[578],seed[66],seed[520],seed[1764],seed[2097],seed[1613],seed[3894],seed[337],seed[3205],seed[3749],seed[628],seed[1395],seed[3222],seed[1409],seed[3680],seed[2340],seed[3986],seed[243],seed[1466],seed[2696],seed[3494],seed[746],seed[1571],seed[1364],seed[2518],seed[2643],seed[378],seed[1401],seed[1667],seed[248],seed[2036],seed[1936],seed[2331],seed[2906],seed[2967],seed[2755],seed[2131],seed[3915],seed[1675],seed[2646],seed[1535],seed[1620],seed[2605],seed[3877],seed[2527],seed[3594],seed[478],seed[3407],seed[1993],seed[1164],seed[484],seed[380],seed[3753],seed[1828],seed[1768],seed[2579],seed[1504],seed[3047],seed[186],seed[1301],seed[3400],seed[2721],seed[563],seed[277],seed[887],seed[1860],seed[1642],seed[3227],seed[3160],seed[1588],seed[1818],seed[4032],seed[3760],seed[3441],seed[1880],seed[528],seed[1943],seed[1458],seed[3751],seed[3702],seed[1067],seed[415],seed[300],seed[2581],seed[2733],seed[2308],seed[1046],seed[3860],seed[466],seed[3114],seed[3598],seed[4023],seed[3945],seed[725],seed[1690],seed[973],seed[1050],seed[2979],seed[502],seed[3352],seed[3308],seed[253],seed[2658],seed[3037],seed[2688],seed[1068],seed[142],seed[3724],seed[3462],seed[133],seed[2497],seed[2731],seed[274],seed[3176],seed[1610],seed[270],seed[392],seed[2935],seed[1702],seed[112],seed[307],seed[1689],seed[2095],seed[1002],seed[1538],seed[1436],seed[156],seed[1810],seed[1157],seed[501],seed[2399],seed[1648],seed[3839],seed[3804],seed[35],seed[1092],seed[554],seed[3310],seed[483],seed[2298],seed[3952],seed[282],seed[3219],seed[331],seed[1908],seed[2730],seed[1583],seed[2005],seed[2788],seed[3049],seed[2145],seed[1753],seed[2100],seed[2986],seed[702],seed[2422],seed[3174],seed[2949],seed[3339],seed[2446],seed[163],seed[3298],seed[2262],seed[1874],seed[3980],seed[3022],seed[3108],seed[2781],seed[1600],seed[3854],seed[757],seed[2743],seed[2342],seed[780],seed[799],seed[1517],seed[4036],seed[926],seed[1482],seed[2933],seed[3563],seed[2182],seed[94],seed[2232],seed[1291],seed[3399],seed[2285],seed[1126],seed[872],seed[2366],seed[1162],seed[1452],seed[824],seed[1240],seed[2580],seed[1379],seed[787],seed[3535],seed[1206],seed[3373],seed[732],seed[3141],seed[1020],seed[1394],seed[3933],seed[1543],seed[3099],seed[933],seed[437],seed[3715],seed[3209],seed[1503],seed[3421],seed[303],seed[3922],seed[2835],seed[3650],seed[3788],seed[386],seed[3490],seed[3082],seed[2374],seed[1565],seed[3743],seed[2663],seed[2426],seed[2598],seed[3165],seed[3414],seed[2913],seed[3552],seed[3549],seed[2983],seed[2396],seed[1983],seed[3542],seed[3102],seed[188],seed[703],seed[717],seed[3427],seed[2457],seed[2459],seed[2700],seed[2136],seed[2744],seed[1055],seed[2453],seed[1998],seed[1418],seed[754],seed[3882],seed[2415],seed[2921],seed[3360],seed[2196],seed[643],seed[2238],seed[822],seed[959],seed[506],seed[438],seed[398],seed[2582],seed[2942],seed[3613],seed[1245],seed[1047],seed[3725],seed[2177],seed[1881],seed[1585],seed[3434],seed[3065],seed[2617],seed[1741],seed[3938],seed[2968],seed[20],seed[920],seed[1801],seed[2498],seed[4072],seed[2657],seed[2263],seed[2635],seed[3005],seed[892],seed[1963],seed[27],seed[4092],seed[516],seed[4013],seed[3169],seed[870],seed[3512],seed[2051],seed[2105],seed[2042],seed[1770],seed[192],seed[1542],seed[2397],seed[1559],seed[421],seed[58],seed[155],seed[3619],seed[2786],seed[2681],seed[2409],seed[3714],seed[219],seed[1172],seed[1121],seed[726],seed[339],seed[2960],seed[919],seed[1557],seed[3217],seed[3772],seed[1918],seed[3832],seed[646],seed[1016],seed[495],seed[982],seed[3491],seed[2260],seed[3392],seed[281],seed[3897],seed[1774],seed[1639],seed[3015],seed[3026],seed[2035],seed[2472],seed[3639],seed[1191],seed[2096],seed[577],seed[217],seed[3446],seed[2085],seed[2784],seed[1520],seed[616],seed[1799],seed[4000],seed[594],seed[1933],seed[1321],seed[2789],seed[2661],seed[448],seed[2545],seed[406],seed[3962],seed[3115],seed[1314],seed[2806],seed[2227],seed[3470],seed[3889],seed[3858],seed[2419],seed[898],seed[2141],seed[1788],seed[1892],seed[738],seed[3155],seed[2412],seed[636],seed[2651],seed[3243],seed[4043],seed[2517],seed[2090],seed[475],seed[1145],seed[917],seed[3793],seed[132],seed[3210],seed[871],seed[709],seed[2286],seed[1477],seed[1851],seed[3323],seed[1045],seed[1579],seed[3762],seed[3572],seed[3106],seed[2938],seed[1723],seed[3687],seed[2269],seed[1666],seed[645],seed[921],seed[1130],seed[3841],seed[195],seed[3095],seed[2275],seed[1578],seed[916],seed[3273],seed[2456],seed[1282],seed[3231],seed[3538],seed[2172],seed[95],seed[1342],seed[663],seed[3701],seed[410],seed[3719],seed[1330],seed[23],seed[1804],seed[811],seed[2574],seed[24],seed[2078],seed[3623],seed[2398],seed[2200],seed[653],seed[739],seed[2296],seed[1814],seed[1064],seed[3211],seed[1512],seed[701],seed[574],seed[1727],seed[113],seed[3990],seed[1400],seed[2793],seed[3982],seed[1817],seed[2108],seed[2951],seed[1439],seed[611],seed[2958],seed[3040],seed[2846],seed[867],seed[2022],seed[1378],seed[3700],seed[1739],seed[3698],seed[2471],seed[3634],seed[1533],seed[2282],seed[239],seed[1805],seed[878],seed[1471],seed[3961],seed[79],seed[2447],seed[593],seed[3705],seed[3953],seed[786],seed[2058],seed[3043],seed[2500],seed[3301],seed[3483],seed[2945],seed[2837],seed[1076],seed[2926],seed[1703],seed[316],seed[3848],seed[3580],seed[3162],seed[497],seed[2102],seed[770],seed[2319],seed[1377],seed[4037],seed[935],seed[1891],seed[265],seed[748],seed[1595],seed[3979],seed[2600],seed[756],seed[3820],seed[3046],seed[1001],seed[1843],seed[2822],seed[474],seed[1144],seed[4046],seed[3194],seed[3935],seed[623],seed[2234],seed[3093],seed[2478],seed[3291],seed[758],seed[2508],seed[1950],seed[4010],seed[2880],seed[1956],seed[52],seed[126],seed[2594],seed[141],seed[1343],seed[3452],seed[913],seed[836],seed[2899],seed[1324],seed[1165],seed[2888],seed[3768],seed[1370],seed[1298],seed[714],seed[4047],seed[1607],seed[3781],seed[981],seed[3058],seed[144],seed[199],seed[2333],seed[1771],seed[1244],seed[2450],seed[3311],seed[1574],seed[2008],seed[2347],seed[3666],seed[4027],seed[2477],seed[1286],seed[3960],seed[2084],seed[3258],seed[2114],seed[3304],seed[678],seed[3557],seed[2692],seed[695],seed[3607],seed[1826],seed[74],seed[2479],seed[2424],seed[2831],seed[2881],seed[433],seed[762],seed[2462],seed[1492],seed[1358],seed[1219],seed[268],seed[3612],seed[706],seed[418],seed[666],seed[2535],seed[114],seed[42],seed[147],seed[2046],seed[3853],seed[1116],seed[3608],seed[581],seed[1671],seed[3419],seed[569],seed[1369],seed[2146],seed[3592],seed[809],seed[216],seed[84],seed[1706],seed[988],seed[661],seed[2709],seed[1732],seed[3364],seed[2233],seed[1832],seed[3268],seed[3034],seed[2386],seed[3396],seed[365],seed[482],seed[1808],seed[3321],seed[583],seed[3097],seed[3477],seed[3502],seed[1457],seed[2395],seed[2],seed[152],seed[1309],seed[1905],seed[2454],seed[1698],seed[1035],seed[1],seed[190],seed[3569],seed[3807],seed[3199],seed[123],seed[3113],seed[2738],seed[202],seed[1118],seed[740],seed[3011],seed[2607],seed[654],seed[672],seed[3653],seed[1320],seed[1778],seed[241],seed[3633],seed[269],seed[1391],seed[1177],seed[2150],seed[470],seed[3277],seed[3378],seed[3823],seed[1949],seed[3849],seed[1955],seed[1563],seed[2727],seed[3312],seed[4071],seed[3754],seed[515],seed[2621],seed[2713],seed[2602],seed[1186],seed[2932],seed[582],seed[254],seed[2593],seed[2373],seed[720],seed[368],seed[2995],seed[3792],seed[4061],seed[3362],seed[1769],seed[2777],seed[496],seed[1684],seed[3548],seed[246],seed[1146],seed[3847],seed[1034],seed[2101],seed[1044],seed[3577],seed[1968],seed[4011],seed[1496],seed[2434],seed[3406],seed[1568],seed[2230],seed[3361],seed[259],seed[845],seed[634],seed[1940],seed[3695],seed[1308],seed[1069],seed[3135],seed[3356],seed[3536],seed[3404],seed[1719],seed[512],seed[257],seed[2192],seed[1700],seed[827],seed[2128],seed[2514],seed[3170],seed[3912],seed[3803],seed[354],seed[1141],seed[1152],seed[3420],seed[3673],seed[1110],seed[1790],seed[320],seed[3934],seed[214],seed[3041],seed[455],seed[1470],seed[3175],seed[641],seed[4015],seed[3503],seed[2247],seed[2293],seed[2082],seed[3787],seed[3487],seed[1926],seed[627],seed[2550],seed[472],seed[3329],seed[1887],seed[1590],seed[2440],seed[764],seed[1674],seed[3726],seed[2390],seed[76],seed[3625],seed[2511],seed[2823],seed[2089],seed[2564],seed[662],seed[3677],seed[2799],seed[831],seed[1350],seed[2666],seed[440],seed[135],seed[3831],seed[603],seed[608],seed[1668],seed[2538],seed[2429],seed[396],seed[2862],seed[3545],seed[2437],seed[93],seed[2253],seed[2917],seed[3507],seed[3439],seed[498],seed[1825],seed[3326],seed[3437],seed[1985],seed[2276],seed[1539],seed[3068],seed[3766],seed[3694],seed[1312],seed[1748],seed[1276],seed[1673],seed[772],seed[1420],seed[1964],seed[2029],seed[41],seed[2798],seed[3266],seed[2155],seed[119],seed[2894],seed[86],seed[304],seed[1904],seed[928],seed[2766],seed[3829],seed[1209],seed[3375],seed[960],seed[4054],seed[3481],seed[2458],seed[1979],seed[1486],seed[3588],seed[3821],seed[2185],seed[2537],seed[2726],seed[3898],seed[733],seed[1082],seed[2569],seed[1709],seed[925],seed[2874],seed[1003],seed[1972],seed[4035],seed[1793],seed[2649],seed[160],seed[103],seed[751],seed[800],seed[1593],seed[915],seed[3458],seed[2436],seed[2869],seed[3193],seed[3879],seed[2838],seed[2092],seed[918],seed[798],seed[3413],seed[951],seed[3863],seed[1975],seed[2417],seed[3264],seed[3045],seed[2499],seed[3624],seed[937],seed[2166],seed[3995],seed[3353],seed[3977],seed[251],seed[346],seed[2118],seed[3746],seed[620],seed[143],seed[2853],seed[3857],seed[2281],seed[127],seed[1037],seed[436],seed[2775],seed[2066],seed[344],seed[1502],seed[3901],seed[2217],seed[1267],seed[2669],seed[366],seed[897],seed[773],seed[2184],seed[2201],seed[2083],seed[3314],seed[1758],seed[3683],seed[3350],seed[1101],seed[3621],seed[26],seed[1526],seed[629],seed[1848],seed[3418],seed[905],seed[1659],seed[1682],seed[2912],seed[2887],seed[399],seed[3246],seed[3916],seed[3524],seed[2769],seed[3275],seed[493],seed[1318],seed[211],seed[1921],seed[3833],seed[2485],seed[213],seed[3496],seed[1188],seed[184],seed[2384],seed[3984],seed[3369],seed[4074],seed[1506],seed[2856],seed[139],seed[461],seed[3657],seed[2064],seed[308],seed[3236],seed[2000],seed[1151],seed[2555],seed[2937],seed[3180],seed[3941],seed[4018],seed[2925],seed[899],seed[1437],seed[1937],seed[3330],seed[680],seed[2294],seed[2024],seed[1902],seed[3454],seed[1000],seed[2616],seed[88],seed[2918],seed[1010],seed[2408],seed[585],seed[3651],seed[335],seed[3381],seed[1767],seed[804],seed[2324],seed[2246],seed[2274],seed[4064],seed[3056],seed[7],seed[1987],seed[2601],seed[3501],seed[3048],seed[2353],seed[1021],seed[3629],seed[3780],seed[1017],seed[4049],seed[2438],seed[499],seed[1977],seed[376],seed[3670],seed[3850],seed[3737],seed[2747],seed[2231],seed[3313],seed[408],seed[1428],seed[1269],seed[1228],seed[3493],seed[2251],seed[2257],seed[1031],seed[3129],seed[2715],seed[1323],seed[2174],seed[3830],seed[173],seed[3796],seed[1519],seed[3061],seed[1265],seed[1839],seed[730],seed[3163],seed[1270],seed[1773],seed[1895],seed[774],seed[2985],seed[2996],seed[4059],seed[271],seed[3927],seed[984],seed[673],seed[2205],seed[1550],seed[1410],seed[468],seed[224],seed[2245],seed[1942],seed[1896],seed[1525],seed[18],seed[3408],seed[955],seed[2543],seed[3985],seed[2159],seed[1742],seed[289],seed[2559],seed[548],seed[2207],seed[785],seed[579],seed[149],seed[3096],seed[1088],seed[2439],seed[3895],seed[968],seed[508],seed[521],seed[2641],seed[1302],seed[2914],seed[3571],seed[3904],seed[3835],seed[2377],seed[3307],seed[1230],seed[1463],seed[3837],seed[3184],seed[3540],seed[3239],seed[1944],seed[503],seed[1441],seed[2833],seed[3606],seed[1147],seed[2520],seed[3125],seed[1432],seed[3260],seed[204],seed[404],seed[1019],seed[2615],seed[1161],seed[2638],seed[1299],seed[3179],seed[299],seed[4038],seed[778],seed[1349],seed[1280],seed[532],seed[4044],seed[1644],seed[264],seed[1416],seed[2026],seed[3654],seed[1782],seed[3968],seed[323],seed[719],seed[82],seed[2198],seed[969],seed[877],seed[207],seed[1934],seed[1930],seed[221],seed[2832],seed[2751],seed[1627],seed[711],seed[3691],seed[4006],seed[340],seed[1890],seed[1665],seed[3116],seed[1140],seed[1057],seed[2972],seed[2506],seed[158],seed[4091],seed[178],seed[2778],seed[2370],seed[2123],seed[1755],seed[2240],seed[3635],seed[1548],seed[3476],seed[4057],seed[614],seed[2599],seed[0],seed[2924],seed[2402],seed[3131],seed[453],seed[130],seed[2783],seed[2327],seed[660],seed[2305],seed[2512],seed[328],seed[302],seed[1204],seed[1852],seed[1919],seed[3672],seed[136],seed[2557],seed[2041],seed[3267],seed[2465],seed[306],seed[745],seed[1408],seed[50],seed[2991],seed[3417],seed[1928],seed[2164],seed[1868],seed[1691],seed[941],seed[3128],seed[2842],seed[3627],seed[1711],seed[1696],seed[2699],seed[3012],seed[454],seed[2705],seed[2801],seed[4069],seed[1053],seed[4030],seed[866],seed[1327],seed[1996],seed[1345],seed[2109],seed[1093],seed[4065],seed[2416],seed[1078],seed[2153],seed[3603],seed[183],seed[4066],seed[2455],seed[1728],seed[1040],seed[3689],seed[353],seed[1091],seed[3252],seed[834],seed[90],seed[3996],seed[954],seed[1952],seed[2040],seed[2065],seed[3038],seed[965],seed[3358],seed[3855],seed[3728],seed[847],seed[3827],seed[696],seed[983],seed[1337],seed[808],seed[3447],seed[1483],seed[1333],seed[3534],seed[1313],seed[3091],seed[2757],seed[2736],seed[2015],seed[3300],seed[617],seed[670],seed[129],seed[3674],seed[3394],seed[3523],seed[1749],seed[389],seed[294],seed[1213],seed[1765],seed[2886],seed[1641],seed[2664],seed[401],seed[881],seed[3468],seed[850],seed[1806],seed[1917],seed[715],seed[3148],seed[3575],seed[2405],seed[2989],seed[458],seed[3218],seed[3000],seed[952],seed[263],seed[551],seed[49],seed[1227],seed[3744],seed[360],seed[637],seed[1498],seed[4014],seed[2662],seed[2139],seed[2909],seed[1351],seed[2577],seed[1406],seed[3002],seed[2898],seed[2704],seed[1969],seed[2361],seed[3690],seed[2915],seed[3325],seed[1072],seed[1203],seed[456],seed[1398],seed[59],seed[3574],seed[3401],seed[324],seed[2488],seed[598],seed[3786],seed[2507],seed[1234],seed[318],seed[633],seed[665],seed[595],seed[325],seed[379],seed[1951],seed[2316],seed[2104],seed[2053],seed[1734],seed[3620],seed[33],seed[3459],seed[1297],seed[3824],seed[349],seed[3931],seed[622],seed[3669],seed[1655],seed[3319],seed[2197],seed[1217],seed[1631],seed[1014],seed[909],seed[1882],seed[2761],seed[3596],seed[4068],seed[167],seed[2750],seed[3112],seed[2191],seed[604],seed[2558],seed[131],seed[319],seed[3771],seed[2977],seed[3188],seed[280],seed[1611],seed[3678],seed[1511],seed[2572],seed[3225],seed[1307],seed[4026],seed[3411],seed[3911],seed[1705],seed[3940],seed[953],seed[1553],seed[2648],seed[1290],seed[227],seed[2335],seed[489],seed[3963],seed[3294],seed[137],seed[2855],seed[89],seed[1685],seed[244],seed[3092],seed[3553],seed[1999],seed[2562],seed[1859],seed[1154],seed[3449],seed[1490],seed[3805],seed[276],seed[220],seed[1075],seed[510],seed[500],seed[2813],seed[3136],seed[1087],seed[2144],seed[3247],seed[1277],seed[1259],seed[2300],seed[2115],seed[3782],seed[1249],seed[707],seed[1124],seed[2765],seed[3430],seed[2267],seed[2608],seed[3685],seed[2866],seed[1194],seed[613],seed[181],seed[3006],seed[2208],seed[326],seed[4052],seed[3903],seed[2423],seed[1266],seed[2759],seed[3366],seed[2032],seed[2536],seed[2264],seed[355],seed[1853],seed[3282],seed[995],seed[361],seed[2461],seed[1854],seed[296],seed[1816],seed[1449],seed[1085],seed[2140],seed[4020],seed[3584],seed[148],seed[1547],seed[1971],seed[1581],seed[2919],seed[1285],seed[3074],seed[2463],seed[460],seed[549],seed[1095],seed[1617],seed[3886],seed[1125],seed[3089],seed[434],seed[1857],seed[2676],seed[2199],seed[1105],seed[1360],seed[1444],seed[1530],seed[1205],seed[1795],seed[1626],seed[3551],seed[4088],seed[3079],seed[3861],seed[2072],seed[3758],seed[397],seed[1923],seed[3717],seed[3951],seed[1293],seed[2425],seed[2007],seed[3457],seed[1056],seed[2540],seed[1893],seed[638],seed[3133],seed[1422],seed[3050],seed[2805],seed[105],seed[2012],seed[943],seed[655],seed[843],seed[1241],seed[708],seed[2711],seed[1243],seed[1913],seed[3713],seed[3943],seed[1558],seed[1182],seed[2844],seed[553],seed[816],seed[1780],seed[3932],seed[2762],seed[2929],seed[3062],seed[3601],seed[3706],seed[3561],seed[2057],seed[2836],seed[226],seed[1621],seed[237],seed[2219],seed[2928],seed[2206],seed[3018],seed[2753],seed[2119],seed[904],seed[3884],seed[1319],seed[3398],seed[2742],seed[741],seed[3819],seed[2796],seed[3518],seed[3759],seed[1138],seed[3974],seed[2586],seed[3573],seed[3384],seed[2722],seed[1763],seed[2381],seed[407],seed[1250],seed[2302],seed[25],seed[1339],seed[1256],seed[1338],seed[1619],seed[3024],seed[3785],seed[2841],seed[2604],seed[1622],seed[54],seed[3206],seed[3259],seed[911],seed[2020],seed[1827],seed[3517],seed[1128],seed[402],seed[367],seed[687],seed[934],seed[2952],seed[1946],seed[3289],seed[3516],seed[3585],seed[1396],seed[2080],seed[2566],seed[2213],seed[2087],seed[3021],seed[2901],seed[2002],seed[3838],seed[1272],seed[3492],seed[768],seed[3320],seed[882],seed[2800],seed[1594],seed[1907],seed[3071],seed[3122],seed[1214],seed[990],seed[3388],seed[3118],seed[1865],seed[3693],seed[3475],seed[3808],seed[2611],seed[3482],seed[1986],seed[3582],seed[1640],seed[3371],seed[3937],seed[3315],seed[4083],seed[3647],seed[667],seed[876],seed[315],seed[2266],seed[1390],seed[2033],seed[755],seed[2625],seed[2130],seed[122],seed[1591],seed[180],seed[3212],seed[2309],seed[3060],seed[596],seed[1454],seed[1570],seed[2549],seed[3905],seed[1080],seed[3004],seed[145],seed[3473],seed[209],seed[2225],seed[3907],seed[403],seed[3716],seed[1796],seed[2418],seed[2167],seed[2341],seed[2045],seed[3656],seed[828],seed[229],seed[1721],seed[2834],seed[795],seed[3667],seed[428],seed[4004],seed[698],seed[2067],seed[75],seed[2226],seed[169],seed[100],seed[3409],seed[3337],seed[1150],seed[1348],seed[3570],seed[2851],seed[519],seed[3727],seed[1381],seed[609],seed[3357],seed[1274],seed[1509],seed[1208],seed[1402],seed[3997],seed[431],seed[657],seed[3098],seed[2328],seed[2810],seed[825],seed[631],seed[118],seed[2103],seed[87],seed[2815],seed[2363],seed[1794],seed[2411],seed[2980],seed[1024],seed[2487],seed[3971],seed[1015],seed[2668],seed[2767],seed[1008],seed[1629],seed[2362],seed[1216],seed[979],seed[2486],seed[597],seed[3547],seed[844],seed[4048],seed[1393],seed[2148],seed[505],seed[1670],seed[936],seed[245],seed[2367],seed[3164],seed[2356],seed[2571],seed[3334],seed[1117],seed[3213],seed[53],seed[2365],seed[3077],seed[3488],seed[2489],seed[647],seed[298],seed[2156],seed[272],seed[3262],seed[3423],seed[3377],seed[2171],seed[1468],seed[3137],seed[3132],seed[2587],seed[1423],seed[3472],seed[1787],seed[1683],seed[2165],seed[345],seed[2371],seed[1676],seed[1582],seed[3117],seed[3834],seed[327],seed[382],seed[2982],seed[3987],seed[3140],seed[2719],seed[3237],seed[1612],seed[417],seed[2680],seed[2435],seed[39],seed[3739],seed[4078],seed[3942],seed[1751],seed[3153],seed[691],seed[846],seed[964],seed[284],seed[2953],seed[1862],seed[2523],seed[200],seed[902],seed[146],seed[2843],seed[3784],seed[601],seed[198],seed[1537],seed[2081],seed[888],seed[1359],seed[526],seed[2242],seed[3899],seed[879],seed[564],seed[818],seed[2858],seed[2152],seed[3280],seed[252],seed[1939],seed[1252],seed[1688],seed[2406],seed[2650],seed[1033],seed[618],seed[3611],seed[2884],seed[1633],seed[2734],seed[4005],seed[36],seed[2277],seed[1103],seed[2613],seed[1435],seed[1442],seed[1296],seed[565],seed[2522],seed[791],seed[1325],seed[2315],seed[863],seed[3978],seed[1647],seed[2444],seed[1462],seed[369],seed[3391],seed[796],seed[793],seed[3478],seed[3800],seed[1635],seed[835],seed[976],seed[1304],seed[3511],seed[171],seed[1586],seed[2687],seed[261],seed[588],seed[3688],seed[1989],seed[1836],seed[3272],seed[523],seed[649],seed[2916],seed[174],seed[961],seed[561],seed[17],seed[3223],seed[78],seed[2821],seed[1238],seed[1136],seed[895],seed[759],seed[2712],seed[2547],seed[2623],seed[4075],seed[1179],seed[749],seed[586],seed[1699],seed[2513],seed[1131],seed[3872],seed[3589],seed[1779],seed[684],seed[560],seed[813],seed[1510],seed[1980],seed[1200],seed[3064],seed[124],seed[729],seed[177],seed[2301],seed[3425],seed[2717],seed[535],seed[3370],seed[416],seed[3506],seed[4007],seed[3017],seed[2748],seed[3202],seed[977],seed[1866],seed[688],seed[3846],seed[752],seed[154],seed[2797],seed[446],seed[3059],seed[2493],seed[2957],seed[893],seed[1375],seed[802],seed[150],seed[765],seed[3382],seed[587],seed[3809],seed[3467],seed[3432],seed[2947],seed[405],seed[2160],seed[639],seed[1176],seed[3293],seed[1809],seed[1160],seed[700],seed[1864],seed[3776],seed[1411],seed[2872],seed[1397],seed[3085],seed[2337],seed[3964],seed[2203],seed[3220],seed[1480],seed[2988],seed[2521],seed[3681],seed[840],seed[1750],seed[1222],seed[3662],seed[1861],seed[2510],seed[1833],seed[3063],seed[2737],seed[2503],seed[1900],seed[3100],seed[2391],seed[2883],seed[1300],seed[632],seed[1807],seed[2178],seed[2376],seed[3198],seed[1499],seed[2678],seed[1746],seed[1005],seed[3692],seed[3271],seed[2708],seed[4062],seed[713],seed[1048],seed[2812],seed[2393],seed[2025],seed[2218],seed[537],seed[1991],seed[3224],seed[2795],seed[2170],seed[414],seed[2466],seed[2496],seed[3887],seed[1210],seed[117],seed[1340],seed[2873],seed[1104],seed[2330],seed[3498],seed[3345],seed[1143],seed[658],seed[3822],seed[4033],seed[1071],seed[3107],seed[3738],seed[333],seed[2934],seed[1284],seed[914],seed[3281],seed[305],seed[4001],seed[3583],seed[838],seed[44],seed[2716],seed[2877],seed[1863],seed[3587],seed[2287],seed[1978],seed[656],seed[681],seed[2970],seed[1198],seed[2318],seed[210],seed[2420],seed[1855],seed[3958],seed[2349],seed[1577],seed[2237],seed[2404],seed[1038],seed[1948],seed[2427],seed[2780],seed[2414],seed[2186],seed[3365],seed[2946],seed[2378],seed[2223],seed[2329],seed[1148],seed[1485],seed[3537],seed[2961],seed[1914],seed[3642],seed[1786],seed[989],seed[1374],seed[3344],seed[1775],seed[1616],seed[3546],seed[383],seed[3124],seed[92],seed[514],seed[1701],seed[373],seed[699],seed[1412],seed[3852],seed[317],seed[3250],seed[884],seed[3504],seed[3296],seed[342],seed[807],seed[3254],seed[1231],seed[2311],seed[3185],seed[1982],seed[3248],seed[3764],seed[2034],seed[3777],seed[2840],seed[357],seed[1306],seed[425],seed[3075],seed[3126],seed[68],seed[1784],seed[1481],seed[1012],seed[2355],seed[3429],seed[3729],seed[2504],seed[1835],seed[689],seed[2074],seed[492],seed[3813],seed[3147],seed[1253],seed[2049],seed[3825],seed[2241],seed[2922],seed[3558],seed[3039],seed[3505],seed[8],seed[2235],seed[1731],seed[4094],seed[3348],seed[2773],seed[1716],seed[3324],seed[2401],seed[3618],seed[1965],seed[3244],seed[2892],seed[2860],seed[96],seed[3461],seed[3568],seed[3665],seed[753],seed[1545],seed[3238],seed[2011],seed[975],seed[3525],seed[1168],seed[419],seed[1058],seed[3908],seed[2895],seed[2261],seed[1598],seed[734],seed[3203],seed[682],seed[2876],seed[949],seed[1247],seed[3615],seed[2467],seed[377],seed[166],seed[3902],seed[3721],seed[1678],seed[1451],seed[1850],seed[2464],seed[3555],seed[1792],seed[2553],seed[1229],seed[225],seed[1041],seed[1812],seed[232],seed[3871],seed[1326],seed[932],seed[1561],seed[297],seed[1341],seed[1007],seed[3870],seed[2820],seed[2694],seed[2997],seed[1677],seed[1514],seed[2243],seed[1139],seed[550],seed[3335],seed[3485],seed[1536],seed[3390],seed[3158],seed[247],seed[2729],seed[2875],seed[1281],seed[3969],seed[939],seed[1417],seed[1988],seed[1687],seed[3207],seed[4021],seed[412],seed[1938],seed[2707],seed[288],seed[473],seed[974],seed[1084],seed[3428],seed[1450],seed[2181],seed[2573],seed[3438],seed[1257],seed[9],seed[31],seed[3867],seed[3290],seed[1329],seed[287],seed[3251],seed[826],seed[829],seed[2891],seed[944],seed[612],seed[889],seed[1884],seed[801],seed[3208],seed[1356],seed[2597],seed[602],seed[1540],seed[222],seed[2289],seed[3649],seed[1875],seed[865],seed[3991],seed[2870],seed[2480],seed[1279],seed[3181],seed[2303],seed[1263],seed[513],seed[3736],seed[3842],seed[423],seed[2852],seed[1941],seed[3906],seed[1576],seed[3696],seed[3609],seed[1883],seed[3981],seed[2673],seed[1730],seed[2516],seed[1844],seed[985],seed[2896],seed[1811],seed[2009],seed[3177],seed[2279],seed[692],seed[1185],seed[3055],seed[2760],seed[2126],seed[504],seed[967],seed[2561],seed[2069],seed[2897],seed[886],seed[3733],seed[2339],seed[3233],seed[3104],seed[3712],seed[29],seed[3463],seed[1066],seed[301],seed[2010],seed[763],seed[2848],seed[1516],seed[3397],seed[1175],seed[1135],seed[3799],seed[1163],seed[2907],seed[3874],seed[1625],seed[1521],seed[862],seed[2332],seed[3235],seed[3495],seed[3878],seed[347],seed[6],seed[2644],seed[1387],seed[63],seed[462],seed[3274],seed[2344],seed[2304],seed[2563],seed[3641],seed[3042],seed[2273],seed[978],seed[2619],seed[3815],seed[1580],seed[3292],seed[2120],seed[3646],seed[4067],seed[3489],seed[3016],seed[4009],seed[3527],seed[1294],seed[3306],seed[571],seed[2674],seed[1011],seed[1223],seed[238],seed[3697],seed[1328],seed[1967],seed[2656],seed[3888],seed[1947],seed[693],seed[1365],seed[894],seed[2849],seed[4073],seed[2050],seed[3305],seed[2505],seed[2578],seed[2596],seed[625],seed[3566],seed[2086],seed[1407],seed[1756],seed[1505],seed[3443],seed[769],seed[273],seed[2830],seed[2244],seed[191],seed[2530],seed[2839],seed[2076],seed[1995],seed[3303],seed[2059],seed[782],seed[3783],seed[3845],seed[3660],seed[710],seed[439],seed[1872],seed[3287],seed[2998],seed[3676],seed[2622],seed[992],seed[3811],seed[1166],seed[3703],seed[1464],seed[2474],seed[3959],seed[875],seed[2077],seed[2603],seed[64],seed[3671],seed[359],seed[3284],seed[2112],seed[285],seed[3288],seed[3790],seed[1260],seed[2252],seed[1858],seed[2070],seed[3031],seed[998],seed[2271],seed[3638],seed[321],seed[947],seed[3166],seed[1924],seed[3054],seed[957],seed[1707],seed[3734],seed[2117],seed[2590],seed[1632],seed[1573],seed[2941],seed[1604],seed[2654],seed[3869],seed[3105],seed[2451],seed[2180],seed[2677],seed[91],seed[1662],seed[2272],seed[48],seed[3216],seed[3032],seed[2359],seed[2375],seed[2056],seed[3893],seed[4070],seed[742],seed[2697],seed[690],seed[3509],seed[2809],seed[2460],seed[1113],seed[2944],seed[3286],seed[3159],seed[1889],seed[573],seed[57],seed[1745],seed[1932],seed[2220],seed[28],seed[2609],seed[589],seed[1424],seed[2690],seed[2037],seed[3090],seed[1115],seed[3775],seed[2048],seed[2653],seed[189],seed[3778],seed[907],seed[3270],seed[2013],seed[1556],seed[1747],seed[2610],seed[4024],seed[4058],seed[3543],seed[443],seed[1661],seed[3909],seed[1086],seed[3081],seed[744],seed[2714],seed[420],seed[1515],seed[2826],seed[1615],seed[712],seed[1193],seed[2254],seed[2640],seed[1567],seed[624],seed[3088],seed[1752],seed[590],seed[2595],seed[1692],seed[2369],seed[3331],seed[1389],seed[2808],seed[1336],seed[3652],seed[3999],seed[948],seed[1489],seed[2211],seed[2016],seed[3632],seed[1802],seed[3789],seed[387],seed[488],seed[4034],seed[34],seed[3631],seed[2556],seed[3072],seed[3828],seed[3600],seed[3617],seed[2321],seed[2133],seed[3966],seed[116],seed[1766],seed[1651],seed[21],seed[3257],seed[1669],seed[1478],seed[3843],seed[3355],seed[4016],seed[206],seed[4019],seed[3151],seed[901],seed[558],seed[3890],seed[2639],seed[3466],seed[619],seed[1376],seed[2222],seed[2728],seed[3559],seed[1030],seed[566],seed[3810],seed[2632],seed[128],seed[336],seed[2554],seed[1736],seed[3057],seed[3892],seed[1974],seed[1465],seed[1733],seed[1431],seed[727],seed[1029],seed[3013],seed[2228],seed[107],seed[1672],seed[4089],seed[2614],seed[2911],seed[4],seed[240],seed[1028],seed[233],seed[2392],seed[803],seed[1901],seed[3992],seed[517],seed[671],seed[790],seed[197],seed[1049],seed[3019],seed[1473],seed[747],seed[987],seed[1929],seed[1899],seed[533],seed[938],seed[2221],seed[559],seed[3033],seed[1623],seed[3709],seed[2268],seed[2132],seed[1710],seed[2068],seed[1953],seed[371],seed[591],seed[3143],seed[3988],seed[3748],seed[1445],seed[3276],seed[1224],seed[555],seed[467],seed[1497],seed[3586],seed[3955],seed[2857],seed[3035],seed[1242],seed[3773],seed[2954],seed[2824],seed[3742],seed[218],seed[3010],seed[2701],seed[2948],seed[1142],seed[2491],seed[922],seed[2627],seed[1114],seed[3581],seed[686],seed[134],seed[3309],seed[3924],seed[839],seed[2749],seed[1712],seed[1054],seed[2670],seed[1127],seed[3918],seed[2183],seed[1523],seed[2179],seed[2325],seed[14],seed[2382],seed[104],seed[1189],seed[669],seed[3186],seed[2740],seed[1822],seed[358],seed[3453],seed[3152],seed[2307],seed[2969],seed[3383],seed[4042],seed[3341],seed[704],seed[2879],seed[1361],seed[1448],seed[3976],seed[694],seed[2278],seed[3970],seed[3679],seed[1597],seed[1158],seed[1460],seed[310],seed[3431],seed[2551],seed[2850],seed[858],seed[394],seed[2043],seed[2389],seed[3230],seed[2667],seed[1572],seed[2388],seed[2482],seed[3003],seed[1475],seed[2920],seed[3684],seed[375],seed[2718],seed[547],seed[2685],seed[2956],seed[606],seed[1658],seed[1903],seed[4003],seed[1992],seed[3150],seed[2091],seed[2413],seed[1871],seed[1879],seed[1686],seed[1488],seed[3261],seed[2671],seed[1120],seed[1781],seed[2620],seed[2476],seed[83],seed[821],seed[2647],seed[760],seed[3479],seed[2368],seed[562],seed[1609],seed[3379],seed[1079],seed[4053],seed[1885],seed[635],seed[1371],seed[2383],seed[390],seed[1199],seed[3655],seed[2116],seed[1190],seed[2149],seed[3747],seed[1036],seed[81],seed[2098],seed[2475],seed[3767],seed[290],seed[1886],seed[72],seed[2019],seed[2939],seed[1419],seed[1443],seed[3295],seed[1346],seed[1645],seed[860],seed[1562],seed[962],seed[3008],seed[1352],seed[923],seed[3658],seed[1415],seed[1211],seed[286],seed[1264],seed[2214],seed[945],seed[1664],seed[463],seed[724],seed[3510],seed[3816],seed[3007],seed[3817],seed[3101],seed[2965],seed[3730],seed[1564],seed[1708],seed[4056],seed[2004],seed[2212],seed[309],seed[370],seed[956],seed[2283],seed[2568],seed[38],seed[1650],seed[3249],seed[3868],seed[1761],seed[1922],seed[737],seed[3593],seed[2930],seed[2284],seed[2993],seed[1382],seed[3067],seed[356],seed[1292],seed[1606],seed[1657],seed[2001],seed[869],seed[3318],seed[2364],seed[1178],seed[910],seed[1427],seed[2215],seed[3440],seed[3084],seed[2421],seed[972],seed[963],seed[2542],seed[1785],seed[1873],seed[2297],seed[2533],seed[3539],seed[2110],seed[2431],seed[3732],seed[2900],seed[3191],seed[2407],seed[3451],seed[1601],seed[777],seed[278],seed[1354],seed[1388],seed[255],seed[3023],seed[441],seed[883],seed[2863],seed[3070],seed[3770],seed[1958],seed[3221],seed[1212],seed[3774],seed[2003],seed[3779],seed[1027],seed[2752],seed[644],seed[3708],seed[820],seed[3],seed[1912],seed[2314],seed[2994],seed[2745],seed[2187],seed[4079],seed[172],seed[4076],seed[1438],seed[575],seed[1099],seed[2682],seed[3178],seed[1106],seed[2163],seed[1528],seed[1959],seed[2306],seed[1221],seed[2758],seed[3722],seed[175],seed[3332],seed[3914],seed[352],seed[931],seed[2176],seed[3550],seed[1976],seed[5],seed[1180],seed[293],seed[2490],seed[4085],seed[761],seed[3387],seed[3336],seed[374],seed[3317],seed[3565],seed[991],seed[2971],seed[797],seed[2675],seed[2062],seed[1119],seed[3359],seed[351],seed[311],seed[2027],seed[3531],seed[640],seed[929],seed[3241],seed[2484],seed[2903],seed[856],seed[3197],seed[3798],seed[1170],seed[2515],seed[2976],seed[1070],seed[3755],seed[1697],seed[1738],seed[650],seed[1009],seed[940],seed[1476],seed[873],seed[1373],seed[1004],seed[1246],seed[1876],seed[3316],seed[542],seed[1815],seed[3349],seed[842],seed[2054],seed[1614],seed[1638],seed[4008],seed[2854],seed[2966],seed[3094],seed[567],seed[43],seed[1403],seed[3499],seed[153],seed[1051],seed[2216],seed[3801],seed[3975],seed[3769],seed[552],seed[3030],seed[3465],seed[3497],seed[735],seed[1605],seed[4039],seed[2882],seed[2531],seed[3422],seed[194],seed[1042],seed[3526],seed[781],seed[3156],seed[2441],seed[2259],seed[1129],seed[1074],seed[3731],seed[3171],seed[1357],seed[851],seed[40],seed[464],seed[2904],seed[1842],seed[69],seed[2137],seed[3412],seed[2867],seed[3145],seed[2018],seed[1453],seed[1271],seed[2352],seed[2771],seed[1023],seed[3599],seed[1869],seed[3110],seed[3025],seed[2168],seed[362],seed[2732],seed[534],seed[2162],seed[2372],seed[3913],seed[1720],seed[3528],seed[1363],seed[442],seed[2779],seed[1910],seed[2483],seed[2878],seed[2470],seed[1355],seed[2552],seed[2962],seed[3297],seed[4060],seed[3604],seed[2134],seed[1159],seed[1233],seed[1646],seed[1513],seed[2343],seed[832],seed[1501],seed[1824],seed[1714],seed[3001],seed[2071],seed[767],seed[903],seed[3930],seed[2589],seed[1426],seed[2079],seed[912],seed[80],seed[3232],seed[3602],seed[3757],seed[291],seed[2583],seed[675],seed[2816],seed[1367],seed[779],seed[3675],seed[1334],seed[201],seed[2358],seed[3484],seed[2725],seed[3643],seed[1331],seed[2693],seed[1153],seed[4080],seed[250],seed[2803],seed[993],seed[1405],seed[4050],seed[3917],seed[106],seed[2794],seed[3965],seed[2313],seed[810],seed[2291],seed[3865],seed[2229],seed[1018],seed[3333],seed[1500],seed[531],seed[2494],seed[3053],seed[2044],seed[599],seed[1945],seed[2636],seed[1220],seed[576],seed[610],seed[970],seed[2905],seed[3947],seed[1994],seed[1743],seed[2819],seed[2585],seed[2859],seed[3134],seed[235],seed[3342],seed[2448],seed[343],seed[4051],seed[182],seed[2129],seed[3130],seed[864],seed[1960],seed[3993],seed[1109],seed[381],seed[1062],seed[3948],seed[479],seed[1332],seed[1507],seed[2239],seed[1800],seed[556],seed[1052],seed[2099],seed[2984],seed[70],seed[4081],seed[2107],seed[422],seed[509],seed[1207],seed[2088],seed[67],seed[60],seed[3957],seed[1587],seed[2628],seed[1421],seed[3157],seed[2990],seed[3616],seed[2868],seed[275],seed[642],seed[1534],seed[3187],seed[3567],seed[3864],seed[1990],seed[1134],seed[450],seed[1544],seed[1715],seed[3532],seed[196],seed[165],seed[11],seed[3253],seed[2385],seed[262],seed[857],seed[2940],seed[2764],seed[447],seed[1618],seed[2400],seed[1275],seed[1628],seed[848],seed[1089],seed[2691],seed[400],seed[522],seed[789],seed[3204],seed[228],seed[999],seed[1925],seed[4087],seed[1554],seed[677],seed[1602],seed[868],seed[110],seed[2710],seed[2927],seed[4022],seed[541],seed[3954],seed[2534],seed[3880],seed[1288],seed[1167],seed[854],seed[384],seed[432],seed[161],seed[3368],seed[1566],seed[1589],seed[1549],seed[545],seed[4084],seed[1372],seed[1195],seed[3245],seed[1834],seed[3229],seed[1202],seed[2502],seed[3578],seed[3424],seed[1729],seed[3876],seed[859],seed[1984],seed[3576],seed[2147],seed[1757],seed[1718],seed[788],seed[3195],seed[3103],seed[4029],seed[2865],seed[1225],seed[2255],seed[3836],seed[1560],seed[242],seed[3127],seed[794],seed[2157],seed[721],seed[986],seed[1909],seed[668],seed[3763],seed[1368],seed[1455],seed[2955],seed[1915],seed[413],seed[570],seed[465],seed[205],seed[108],seed[2312],seed[2169],seed[3146],seed[2346],seed[350],seed[2686],seed[1694],seed[511],seed[363],seed[332],seed[2014],seed[2061],seed[3707],seed[223],seed[1201],seed[3562],seed[1073],seed[230],seed[1303],seed[3340],seed[1232],seed[1107],seed[61],seed[2121],seed[891],seed[3885],seed[1278],seed[3925],seed[3009],seed[3640],seed[1713],seed[728],seed[3896],seed[121],seed[322],seed[3167],seed[3234],seed[792],seed[830],seed[1108],seed[3520],seed[236],seed[3862],seed[2814],seed[805],seed[2250],seed[2629],seed[2449],seed[722],seed[3926],seed[2576],seed[2151],seed[783],seed[176],seed[330],seed[258],seed[2790],seed[1803],seed[2908],seed[1289],seed[1187],seed[3756],seed[3590],seed[1935],seed[1762],seed[3405],seed[1096],seed[4002],seed[705],seed[2588],seed[157],seed[1760],seed[3078],seed[3374],seed[4082],seed[385],seed[3471],seed[718],seed[3591],seed[2665],seed[2338],seed[2964],seed[607],seed[430],seed[2584],seed[1174],seed[3797],seed[2073],seed[1173],seed[2999],seed[2931],seed[4095],seed[659],seed[557],seed[19],seed[1484],seed[1603],seed[3508],seed[2357],seed[592],seed[815],seed[231],seed[885],seed[2861],seed[1215],seed[3069],seed[1392],seed[580],seed[3723],seed[3844],seed[2236],seed[1634],seed[338],seed[2811],seed[1261],seed[3279],seed[2360],seed[3989],seed[2548],seed[1552],seed[2322],seed[2936],seed[3051],seed[1060],seed[477],seed[2893],seed[1798],seed[3283],seed[2060],seed[4063],seed[648],seed[861],seed[2154],seed[2817],seed[2143],seed[2943],seed[334],seed[544],seed[743],seed[1663],seed[2890],seed[3172],seed[1097],seed[1032],seed[2351],seed[853],seed[1446],seed[279],seed[1831],seed[1636],seed[817],seed[716],seed[2209],seed[1006],seed[65],seed[2354],seed[2791],seed[2787],seed[2756],seed[2094],seed[3610],seed[4028],seed[16],seed[85],seed[2889],seed[819],seed[1273],seed[1433],seed[1653],seed[3087],seed[3818],seed[849],seed[1656],seed[292],seed[3474],seed[1897],seed[2442],seed[1740],seed[1043],seed[2299],seed[459],seed[1171],seed[2776],seed[1239],seed[1414],seed[1981],seed[451],seed[56],seed[2288],seed[3189],seed[3020],seed[4077],seed[1777],seed[2075],seed[3950],seed[1474],seed[1970],seed[45],seed[2720],seed[1316],seed[3385],seed[2804],seed[775],seed[584],seed[185],seed[2224],seed[162],seed[2735],seed[3367],seed[1380],seed[3735],seed[481],seed[2871],seed[4031],seed[2702],seed[2978],seed[3302],seed[3791],seed[3579],seed[2524],seed[3663],seed[3111],seed[2334],seed[98],seed[2541],seed[2975],seed[771],seed[3664],seed[1100],seed[1584],seed[1830],seed[1823],seed[3190],seed[1957],seed[1819],seed[3347],seed[3605],seed[3873],seed[2741],seed[2612],seed[2492],seed[1704],seed[546],seed[3998],seed[1624],seed[723],seed[3029],seed[3856],seed[3944],seed[51],seed[1531],seed[766],seed[2950],seed[212],seed[187],seed[1112],seed[3444],seed[449],seed[996],seed[3802],seed[3327],seed[2093],seed[2973],seed[256],seed[1888],seed[2345],seed[3752],seed[312],seed[3946],seed[1181],seed[3480],seed[1493],seed[2724],seed[3564],seed[2672],seed[1467],seed[615],seed[3704],seed[529],seed[1637],seed[1254],seed[2193],seed[3415],seed[3044],seed[2630],seed[2626],seed[1838],seed[1846],seed[3628],seed[3120]}),
        .cross_prob(cross_prob),
        .codeword(codeword7),
        .received(received7)
        );
        
    bsc bsc8(
        .clk(clk),
        .reset(reset),
        .seed({seed[2128],seed[2719],seed[1599],seed[3598],seed[1369],seed[1503],seed[1622],seed[241],seed[2621],seed[1680],seed[2037],seed[3670],seed[3210],seed[3434],seed[3846],seed[22],seed[3829],seed[2936],seed[2283],seed[1910],seed[1088],seed[3817],seed[462],seed[3080],seed[1689],seed[3419],seed[150],seed[1999],seed[273],seed[957],seed[3488],seed[1798],seed[1460],seed[3892],seed[1277],seed[3740],seed[2261],seed[3403],seed[2206],seed[1959],seed[255],seed[2183],seed[504],seed[3681],seed[2625],seed[2184],seed[3145],seed[1579],seed[3156],seed[3855],seed[2990],seed[2319],seed[2314],seed[2321],seed[4081],seed[3966],seed[1373],seed[1051],seed[2536],seed[2058],seed[2520],seed[989],seed[2696],seed[3352],seed[565],seed[92],seed[3591],seed[2138],seed[2063],seed[2578],seed[1748],seed[1279],seed[956],seed[60],seed[3884],seed[2948],seed[2142],seed[1254],seed[1833],seed[455],seed[2710],seed[2714],seed[2753],seed[1333],seed[1349],seed[2407],seed[1614],seed[2020],seed[1233],seed[3602],seed[2734],seed[550],seed[1451],seed[673],seed[4058],seed[1228],seed[2120],seed[1640],seed[3933],seed[2046],seed[1057],seed[3465],seed[2608],seed[2829],seed[18],seed[1371],seed[3249],seed[1558],seed[2452],seed[3706],seed[1027],seed[703],seed[1884],seed[269],seed[864],seed[2295],seed[2551],seed[3504],seed[2950],seed[441],seed[2945],seed[2332],seed[927],seed[2777],seed[2679],seed[2790],seed[928],seed[3556],seed[2723],seed[2126],seed[3848],seed[1975],seed[1453],seed[1791],seed[1545],seed[6],seed[1583],seed[171],seed[2351],seed[2820],seed[522],seed[1463],seed[1977],seed[1040],seed[3734],seed[3317],seed[2812],seed[3111],seed[1025],seed[1500],seed[373],seed[1416],seed[3195],seed[2534],seed[629],seed[606],seed[1817],seed[3801],seed[1571],seed[595],seed[2703],seed[839],seed[3028],seed[2430],seed[1075],seed[562],seed[1466],seed[3522],seed[238],seed[1816],seed[614],seed[915],seed[2403],seed[2983],seed[2417],seed[2739],seed[648],seed[110],seed[2494],seed[2080],seed[714],seed[2911],seed[2055],seed[712],seed[2047],seed[807],seed[3297],seed[3222],seed[936],seed[1178],seed[3004],seed[1395],seed[3753],seed[3112],seed[157],seed[3253],seed[1449],seed[2666],seed[1674],seed[2081],seed[878],seed[95],seed[2862],seed[1273],seed[615],seed[3225],seed[2641],seed[1157],seed[1991],seed[530],seed[2467],seed[2928],seed[2560],seed[2962],seed[2176],seed[3068],seed[676],seed[747],seed[3362],seed[474],seed[3940],seed[2994],seed[63],seed[3359],seed[2043],seed[66],seed[534],seed[3217],seed[2012],seed[1208],seed[1313],seed[2432],seed[2297],seed[3197],seed[651],seed[729],seed[1870],seed[459],seed[374],seed[3491],seed[1468],seed[2339],seed[3011],seed[1754],seed[3533],seed[457],seed[2672],seed[1341],seed[781],seed[3354],seed[780],seed[2459],seed[1276],seed[3127],seed[3313],seed[632],seed[3766],seed[853],seed[206],seed[2762],seed[1873],seed[1655],seed[963],seed[2463],seed[2511],seed[718],seed[2033],seed[1865],seed[896],seed[4084],seed[851],seed[1549],seed[1302],seed[3094],seed[608],seed[2294],seed[1159],seed[3452],seed[2499],seed[3511],seed[1670],seed[3315],seed[1268],seed[342],seed[1255],seed[3535],seed[3121],seed[563],seed[997],seed[738],seed[2262],seed[1400],seed[1196],seed[3496],seed[200],seed[210],seed[3660],seed[3852],seed[2298],seed[2835],seed[1770],seed[1906],seed[2858],seed[419],seed[3264],seed[2588],seed[3270],seed[477],seed[2250],seed[1952],seed[3189],seed[3229],seed[1695],seed[1829],seed[3258],seed[3320],seed[452],seed[14],seed[978],seed[222],seed[2445],seed[3446],seed[918],seed[1516],seed[3685],seed[672],seed[3795],seed[2690],seed[3974],seed[2854],seed[3097],seed[188],seed[1652],seed[1024],seed[3584],seed[964],seed[285],seed[1650],seed[1984],seed[1712],seed[2747],seed[1121],seed[2875],seed[3478],seed[1942],seed[2242],seed[1493],seed[3782],seed[2389],seed[2521],seed[971],seed[2076],seed[488],seed[3269],seed[952],seed[3894],seed[2497],seed[1948],seed[2068],seed[2609],seed[3891],seed[3783],seed[3861],seed[3585],seed[3199],seed[2617],seed[2161],seed[2356],seed[1734],seed[2164],seed[4072],seed[253],seed[824],seed[2519],seed[600],seed[3445],seed[3272],seed[2042],seed[503],seed[3730],seed[443],seed[4085],seed[3343],seed[3404],seed[1735],seed[3221],seed[3798],seed[3560],seed[3658],seed[47],seed[903],seed[2373],seed[2999],seed[2611],seed[857],seed[3486],seed[1348],seed[3167],seed[3615],seed[3530],seed[2400],seed[1342],seed[558],seed[3365],seed[2248],seed[3529],seed[838],seed[3400],seed[435],seed[3880],seed[3295],seed[2132],seed[1358],seed[3960],seed[4022],seed[2985],seed[3757],seed[763],seed[2901],seed[1499],seed[2638],seed[2343],seed[2992],seed[1198],seed[3071],seed[65],seed[2119],seed[256],seed[2268],seed[646],seed[1308],seed[1144],seed[2558],seed[3661],seed[3752],seed[340],seed[931],seed[771],seed[2549],seed[106],seed[4054],seed[2413],seed[2310],seed[1298],seed[3555],seed[1262],seed[1737],seed[3634],seed[1047],seed[2289],seed[3517],seed[1114],seed[1854],seed[80],seed[634],seed[2867],seed[846],seed[3649],seed[766],seed[3561],seed[3854],seed[3025],seed[3012],seed[3727],seed[2073],seed[658],seed[3509],seed[3628],seed[2731],seed[3886],seed[2853],seed[2898],seed[299],seed[2648],seed[752],seed[1464],seed[3169],seed[3218],seed[1710],seed[1322],seed[29],seed[4042],seed[1123],seed[3970],seed[368],seed[3984],seed[2504],seed[756],seed[3226],seed[1885],seed[2473],seed[1469],seed[298],seed[2141],seed[2576],seed[3856],seed[553],seed[1133],seed[580],seed[1393],seed[3659],seed[3613],seed[3168],seed[2088],seed[4094],seed[3000],seed[1370],seed[1146],seed[751],seed[2290],seed[3402],seed[152],seed[26],seed[2426],seed[3729],seed[2282],seed[1796],seed[3116],seed[707],seed[2158],seed[1623],seed[1925],seed[3069],seed[3041],seed[3441],seed[2972],seed[2626],seed[3709],seed[3472],seed[1647],seed[1437],seed[2779],seed[1904],seed[3914],seed[906],seed[105],seed[333],seed[3952],seed[3991],seed[2360],seed[3859],seed[1544],seed[955],seed[736],seed[3497],seed[1245],seed[1264],seed[55],seed[1244],seed[576],seed[4089],seed[2085],seed[2701],seed[1964],seed[381],seed[427],seed[3677],seed[1908],seed[1278],seed[3583],seed[1092],seed[2124],seed[3484],seed[190],seed[2107],seed[2181],seed[2932],seed[863],seed[2730],seed[2514],seed[1174],seed[3463],seed[2218],seed[557],seed[1926],seed[4032],seed[3487],seed[885],seed[3872],seed[3995],seed[120],seed[2197],seed[3640],seed[2361],seed[231],seed[2450],seed[1768],seed[3345],seed[509],seed[2897],seed[4091],seed[620],seed[19],seed[297],seed[1501],seed[631],seed[996],seed[1922],seed[117],seed[2386],seed[1741],seed[2584],seed[3067],seed[1588],seed[2196],seed[1830],seed[2515],seed[2154],seed[1511],seed[2293],seed[3701],seed[3245],seed[3899],seed[900],seed[2996],seed[2675],seed[2964],seed[1211],seed[1147],seed[1087],seed[2163],seed[2175],seed[3163],seed[1913],seed[3302],seed[1131],seed[3896],seed[539],seed[679],seed[3776],seed[1386],seed[2900],seed[486],seed[2031],seed[1136],seed[2030],seed[2751],seed[3347],seed[216],seed[4050],seed[1299],seed[2995],seed[3637],seed[2337],seed[146],seed[2772],seed[103],seed[3526],seed[1574],seed[929],seed[3616],seed[3483],seed[3394],seed[2442],seed[1895],seed[2843],seed[827],seed[335],seed[3085],seed[2891],seed[148],seed[1746],seed[1852],seed[1832],seed[3372],seed[1941],seed[1072],seed[1484],seed[1070],seed[1568],seed[3066],seed[652],seed[1032],seed[841],seed[3608],seed[1801],seed[882],seed[1241],seed[1195],seed[1855],seed[1965],seed[3550],seed[3905],seed[2698],seed[362],seed[2699],seed[2317],seed[1170],seed[3287],seed[1557],seed[3206],seed[1728],seed[3519],seed[3430],seed[1532],seed[2465],seed[3309],seed[828],seed[3883],seed[3840],seed[1792],seed[487],seed[516],seed[165],seed[2899],seed[2967],seed[3948],seed[3170],seed[1073],seed[2629],seed[2251],seed[13],seed[2802],seed[2688],seed[607],seed[689],seed[1939],seed[949],seed[659],seed[3024],seed[1316],seed[1985],seed[999],seed[811],seed[4071],seed[2870],seed[350],seed[782],seed[423],seed[2712],seed[1398],seed[3062],seed[496],seed[1200],seed[69],seed[2436],seed[3393],seed[3339],seed[149],seed[965],seed[3209],seed[1215],seed[531],seed[3275],seed[3676],seed[1867],seed[586],seed[3621],seed[1857],seed[674],seed[2968],seed[1766],seed[2487],seed[3668],seed[945],seed[1573],seed[1366],seed[2502],seed[4045],seed[3707],seed[1793],seed[1292],seed[3458],seed[476],seed[3420],seed[2764],seed[1809],seed[2949],seed[988],seed[1296],seed[2903],seed[1321],seed[1183],seed[3188],seed[3379],seed[1699],seed[2257],seed[761],seed[193],seed[1752],seed[1896],seed[2274],seed[191],seed[3983],seed[3841],seed[283],seed[1848],seed[1745],seed[1052],seed[861],seed[2344],seed[3325],seed[732],seed[2071],seed[139],seed[1150],seed[3645],seed[3134],seed[425],seed[3811],seed[1633],seed[2002],seed[995],seed[2976],seed[795],seed[3579],seed[2546],seed[874],seed[182],seed[3407],seed[3712],seed[2615],seed[3527],seed[3408],seed[624],seed[3010],seed[2633],seed[623],seed[1161],seed[2346],seed[2890],seed[301],seed[1894],seed[1345],seed[426],seed[3459],seed[410],seed[2434],seed[1335],seed[3279],seed[1225],seed[2785],seed[643],seed[3961],seed[2823],seed[3946],seed[3182],seed[2482],seed[2377],seed[2309],seed[3962],seed[3166],seed[3026],seed[3557],seed[2709],seed[681],seed[1109],seed[1141],seed[2050],seed[726],seed[2708],seed[3719],seed[1337],seed[2622],seed[1617],seed[3630],seed[167],seed[1664],seed[33],seed[3351],seed[1062],seed[3745],seed[511],seed[3830],seed[3457],seed[2736],seed[1424],seed[1928],seed[1387],seed[324],seed[1786],seed[1272],seed[2117],seed[3323],seed[2249],seed[3534],seed[2906],seed[1003],seed[2078],seed[3439],seed[2077],seed[2643],seed[3870],seed[168],seed[3687],seed[237],seed[992],seed[4002],seed[1654],seed[1325],seed[589],seed[1307],seed[2475],seed[3185],seed[2391],seed[2657],seed[205],seed[2004],seed[3796],seed[3043],seed[3036],seed[1392],seed[1478],seed[1740],seed[556],seed[1524],seed[847],seed[3626],seed[2902],seed[1899],seed[2563],seed[3399],seed[404],seed[246],seed[3818],seed[3409],seed[3376],seed[1651],seed[3747],seed[71],seed[1555],seed[1911],seed[1760],seed[282],seed[719],seed[3921],seed[454],seed[1600],seed[3479],seed[341],seed[264],seed[258],seed[1982],seed[2203],seed[3032],seed[3001],seed[1045],seed[3710],seed[602],seed[2061],seed[2583],seed[2474],seed[3777],seed[3629],seed[2864],seed[533],seed[1636],seed[2811],seed[135],seed[2469],seed[926],seed[891],seed[1730],seed[2654],seed[378],seed[2569],seed[1005],seed[1056],seed[3361],seed[1021],seed[123],seed[275],seed[88],seed[2205],seed[3528],seed[1738],seed[2828],seed[3773],seed[987],seed[555],seed[639],seed[1759],seed[3797],seed[4065],seed[3341],seed[3505],seed[1627],seed[2941],seed[3332],seed[1637],seed[981],seed[2522],seed[2246],seed[609],seed[116],seed[1667],seed[1990],seed[3378],seed[2086],seed[1465],seed[3215],seed[1621],seed[1969],seed[2800],seed[2926],seed[1630],seed[2750],seed[2732],seed[2610],seed[3122],seed[377],seed[2278],seed[2340],seed[3271],seed[1490],seed[3058],seed[3577],seed[1135],seed[384],seed[2997],seed[3383],seed[2122],seed[3037],seed[1715],seed[3609],seed[3057],seed[3211],seed[2632],seed[1180],seed[3778],seed[1285],seed[2481],seed[1175],seed[3240],seed[4008],seed[85],seed[1860],seed[1962],seed[1641],seed[3410],seed[3698],seed[3280],seed[3002],seed[3562],seed[1644],seed[2943],seed[2462],seed[471],seed[585],seed[2556],seed[3614],seed[107],seed[2861],seed[1696],seed[1560],seed[2669],seed[2496],seed[352],seed[1596],seed[2880],seed[1584],seed[4043],seed[1129],seed[2857],seed[393],seed[3329],seed[1878],seed[597],seed[2051],seed[1126],seed[1886],seed[3088],seed[3089],seed[2108],seed[1826],seed[2946],seed[2005],seed[2774],seed[1811],seed[2001],seed[2939],seed[1638],seed[2191],seed[173],seed[1328],seed[875],seed[913],seed[2815],seed[749],seed[1933],seed[3131],seed[3101],seed[1818],seed[3785],seed[2984],seed[178],seed[1893],seed[1054],seed[1412],seed[445],seed[3741],seed[490],seed[3391],seed[3267],seed[217],seed[37],seed[3784],seed[1429],seed[2630],seed[4049],seed[1679],seed[230],seed[1601],seed[1267],seed[2238],seed[3780],seed[3909],seed[2171],seed[3114],seed[1452],seed[2507],seed[3596],seed[3824],seed[3823],seed[1678],seed[227],seed[28],seed[3652],seed[3423],seed[2613],seed[166],seed[2908],seed[1749],seed[2553],seed[3429],seed[572],seed[3130],seed[3033],seed[344],seed[1001],seed[1079],seed[1782],seed[3319],seed[3930],seed[1502],seed[3969],seed[2003],seed[2415],seed[2026],seed[1781],seed[627],seed[1026],seed[3646],seed[656],seed[3009],seed[1360],seed[3413],seed[541],seed[3926],seed[1645],seed[2069],seed[2328],seed[197],seed[2451],seed[3139],seed[2577],seed[3839],seed[2098],seed[1937],seed[2279],seed[1838],seed[1890],seed[938],seed[723],seed[3832],seed[787],seed[3427],seed[429],seed[4056],seed[912],seed[1237],seed[1098],seed[919],seed[954],seed[3181],seed[1841],seed[3187],seed[3506],seed[2850],seed[1763],seed[785],seed[3672],seed[3330],seed[2199],seed[1872],seed[2683],seed[2148],seed[794],seed[1102],seed[1534],seed[2215],seed[3688],seed[1018],seed[768],seed[1739],seed[3768],seed[1543],seed[300],seed[1000],seed[3897],seed[1779],seed[3428],seed[3165],seed[3695],seed[969],seed[2682],seed[3788],seed[3931],seed[4063],seed[986],seed[1954],seed[692],seed[3406],seed[3553],seed[3549],seed[1971],seed[1869],seed[917],seed[3792],seed[402],seed[1577],seed[1293],seed[2716],seed[367],seed[933],seed[665],seed[372],seed[1023],seed[2580],seed[3142],seed[1955],seed[4090],seed[343],seed[1152],seed[2485],seed[3495],seed[1720],seed[1592],seed[1140],seed[2168],seed[3989],seed[3806],seed[1431],seed[748],seed[2054],seed[1874],seed[1363],seed[2027],seed[543],seed[3851],seed[305],seed[3543],seed[83],seed[3597],seed[3091],seed[2425],seed[3665],seed[3431],seed[770],seed[1067],seed[2678],seed[1918],seed[3308],seed[2363],seed[1414],seed[4016],seed[3135],seed[104],seed[2844],seed[1265],seed[1691],seed[4014],seed[3070],seed[2492],seed[1483],seed[3935],seed[3760],seed[3019],seed[2767],seed[3641],seed[391],seed[2052],seed[3433],seed[3518],seed[3369],seed[1488],seed[357],seed[2631],seed[2149],seed[1665],seed[1317],seed[2285],seed[428],seed[3230],seed[3751],seed[760],seed[813],seed[3054],seed[240],seed[2303],seed[2754],seed[127],seed[112],seed[1344],seed[169],seed[1350],seed[549],seed[223],seed[271],seed[3395],seed[2595],seed[409],seed[3900],seed[2667],seed[2889],seed[662],seed[1275],seed[2572],seed[2190],seed[2133],seed[4093],seed[304],seed[613],seed[626],seed[1716],seed[3455],seed[3490],seed[1286],seed[2784],seed[517],seed[2973],seed[2495],seed[592],seed[3076],seed[2048],seed[2449],seed[1381],seed[3539],seed[848],seed[126],seed[3732],seed[2049],seed[1297],seed[1615],seed[3387],seed[1987],seed[1356],seed[705],seed[3653],seed[411],seed[1772],seed[61],seed[1230],seed[2437],seed[3034],seed[2381],seed[582],seed[1154],seed[128],seed[2816],seed[2269],seed[3064],seed[3655],seed[3086],seed[243],seed[2130],seed[336],seed[311],seed[618],seed[1042],seed[3889],seed[1940],seed[2228],seed[1821],seed[158],seed[2292],seed[1034],seed[1718],seed[3177],seed[2471],seed[856],seed[1055],seed[849],seed[2618],seed[2466],seed[2333],seed[279],seed[115],seed[973],seed[96],seed[3631],seed[1082],seed[3128],seed[880],seed[3467],seed[3397],seed[1213],seed[265],seed[3620],seed[1132],seed[650],seed[1086],seed[2147],seed[561],seed[2349],seed[291],seed[1572],seed[2684],seed[3713],seed[347],seed[2256],seed[1970],seed[1492],seed[3237],seed[817],seed[2813],seed[2888],seed[4035],seed[194],seed[2134],seed[327],seed[3462],seed[1866],seed[2272],seed[3642],seed[2179],seed[1404],seed[3243],seed[1256],seed[1812],seed[1188],seed[2725],seed[2390],seed[3794],seed[1435],seed[2804],seed[907],seed[184],seed[734],seed[1015],seed[3007],seed[2752],seed[3865],seed[1112],seed[3636],seed[3375],seed[2411],seed[461],seed[1145],seed[2165],seed[1642],seed[3567],seed[2029],seed[1331],seed[2245],seed[943],seed[4067],seed[3384],seed[1074],seed[2484],seed[3647],seed[108],seed[1871],seed[2616],seed[3589],seed[1512],seed[3895],seed[2221],seed[2925],seed[437],seed[3702],seed[2554],seed[2423],seed[3761],seed[1708],seed[3077],seed[4051],seed[2393],seed[737],seed[2448],seed[1729],seed[358],seed[1656],seed[379],seed[2776],seed[3986],seed[2345],seed[491],seed[1515],seed[2498],seed[953],seed[2532],seed[3083],seed[3913],seed[829],seed[524],seed[2733],seed[3749],seed[3575],seed[1542],seed[2186],seed[1011],seed[823],seed[1936],seed[2100],seed[3881],seed[2302],seed[1427],seed[1261],seed[453],seed[4001],seed[185],seed[960],seed[830],seed[1007],seed[741],seed[189],seed[415],seed[1269],seed[17],seed[254],seed[434],seed[1081],seed[1802],seed[1326],seed[442],seed[67],seed[2311],seed[2072],seed[1458],seed[2860],seed[1059],seed[1593],seed[2022],seed[833],seed[1446],seed[444],seed[2605],seed[1517],seed[212],seed[1038],seed[3079],seed[3153],seed[1153],seed[3968],seed[3787],seed[2674],seed[4],seed[1433],seed[288],seed[276],seed[3065],seed[1657],seed[1457],seed[909],seed[2797],seed[869],seed[406],seed[3082],seed[1439],seed[2483],seed[2905],seed[337],seed[225],seed[1823],seed[3039],seed[968],seed[816],seed[2472],seed[201],seed[1362],seed[3255],seed[1138],seed[2307],seed[696],seed[302],seed[1496],seed[717],seed[1778],seed[2722],seed[1530],seed[2713],seed[90],seed[3835],seed[686],seed[1916],seed[3965],seed[515],seed[2952],seed[1947],seed[868],seed[1085],seed[176],seed[3893],seed[3678],seed[3492],seed[750],seed[1595],seed[1807],seed[3820],seed[1380],seed[2944],seed[1221],seed[722],seed[4088],seed[53],seed[2718],seed[403],seed[560],seed[4044],seed[1078],seed[1019],seed[2461],seed[860],seed[1020],seed[3838],seed[892],seed[2136],seed[1388],seed[1727],seed[3277],seed[680],seed[2229],seed[2527],seed[500],seed[1039],seed[2545],seed[1960],seed[1538],seed[1634],seed[2167],seed[2503],seed[1181],seed[1725],seed[1139],seed[2661],seed[2145],seed[1688],seed[1201],seed[1546],seed[3117],seed[2934],seed[2429],seed[3759],seed[3016],seed[3172],seed[759],seed[3418],seed[685],seed[2300],seed[2094],seed[1923],seed[3074],seed[2839],seed[187],seed[859],seed[902],seed[805],seed[3417],seed[1455],seed[3919],seed[2446],seed[3541],seed[3502],seed[1049],seed[3202],seed[1723],seed[2101],seed[3132],seed[1119],seed[2988],seed[1474],seed[130],seed[2574],seed[2548],seed[2991],seed[611],seed[35],seed[972],seed[835],seed[3592],seed[2367],seed[48],seed[1158],seed[3224],seed[1162],seed[2066],seed[1258],seed[2827],seed[3936],seed[3618],seed[2110],seed[2517],seed[1755],seed[2539],seed[3885],seed[3364],seed[4046],seed[2371],seed[1002],seed[2477],seed[3873],seed[3573],seed[3042],seed[2277],seed[2612],seed[2280],seed[3736],seed[3092],seed[837],seed[4070],seed[2916],seed[2918],seed[3355],seed[2960],seed[366],seed[2129],seed[744],seed[3610],seed[2045],seed[588],seed[3363],seed[1312],seed[2213],seed[1339],seed[4020],seed[3254],seed[3027],seed[351],seed[1988],seed[2938],seed[1184],seed[3571],seed[2506],seed[1359],seed[2571],seed[1620],seed[2304],seed[2422],seed[363],seed[3450],seed[3476],seed[521],seed[2881],seed[2769],seed[776],seed[1856],seed[75],seed[767],seed[2935],seed[274],seed[1064],seed[1619],seed[2464],seed[1639],seed[125],seed[2872],seed[1476],seed[1974],seed[3971],seed[2760],seed[826],seed[289],seed[1846],seed[1762],seed[697],seed[803],seed[1669],seed[801],seed[345],seed[3808],seed[3774],seed[1677],seed[2805],seed[2338],seed[3356],seed[1521],seed[2636],seed[1949],seed[3102],seed[644],seed[2399],seed[1352],seed[323],seed[3120],seed[3673],seed[3699],seed[2385],seed[2624],seed[1487],seed[209],seed[1649],seed[3198],seed[3358],seed[1330],seed[2755],seed[4003],seed[598],seed[481],seed[2222],seed[1525],seed[3957],seed[2707],seed[1514],seed[4005],seed[1683],seed[2234],seed[2267],seed[731],seed[3157],seed[3105],seed[671],seed[3876],seed[1858],seed[181],seed[1658],seed[552],seed[3680],seed[2143],seed[3396],seed[655],seed[2808],seed[4057],seed[3008],seed[1430],seed[1950],seed[180],seed[786],seed[450],seed[2884],seed[260],seed[2728],seed[1413],seed[706],seed[2187],seed[2146],seed[499],seed[1409],seed[1438],seed[316],seed[1410],seed[3314],seed[2288],seed[1014],seed[1378],seed[3412],seed[1205],seed[1220],seed[204],seed[1450],seed[3328],seed[4095],seed[2478],seed[98],seed[1897],seed[2324],seed[473],seed[2153],seed[2336],seed[2568],seed[2526],seed[3906],seed[3246],seed[3178],seed[3624],seed[1537],seed[3866],seed[420],seed[3836],seed[1217],seed[4073],seed[1721],seed[3180],seed[538],seed[3235],seed[3371],seed[3090],seed[3878],seed[2118],seed[49],seed[3453],seed[1567],seed[2264],seed[3104],seed[1690],seed[2253],seed[495],seed[3635],seed[3879],seed[3548],seed[3063],seed[1029],seed[1847],seed[1605],seed[1709],seed[510],seed[2543],seed[742],seed[2642],seed[2489],seed[1840],seed[2299],seed[975],seed[2123],seed[2695],seed[3435],seed[603],seed[3800],seed[799],seed[698],seed[1461],seed[3093],seed[2687],seed[1612],seed[3939],seed[1684],seed[3059],seed[396],seed[4077],seed[1570],seed[2470],seed[3190],seed[383],seed[2192],seed[1017],seed[2057],seed[1836],seed[2789],seed[244],seed[3993],seed[2216],seed[3331],seed[2570],seed[174],seed[1790],seed[3964],seed[2676],seed[2510],seed[3918],seed[1240],seed[2034],seed[1518],seed[2693],seed[3547],seed[2178],seed[380],seed[2064],seed[3607],seed[898],seed[4087],seed[2301],seed[2263],seed[77],seed[962],seed[548],seed[1536],seed[2270],seed[1475],seed[431],seed[1309],seed[4011],seed[1310],seed[132],seed[1602],seed[2056],seed[529],seed[4017],seed[1130],seed[1685],seed[3718],seed[4026],seed[1613],seed[1459],seed[3988],seed[3151],seed[3942],seed[3256],seed[3985],seed[2023],seed[2070],seed[1610],seed[502],seed[1726],seed[4021],seed[1374],seed[3941],seed[467],seed[1440],seed[3155],seed[56],seed[2041],seed[3531],seed[3040],seed[940],seed[1243],seed[4025],seed[242],seed[1785],seed[3587],seed[1861],seed[2160],seed[2308],seed[2018],seed[3693],seed[1473],seed[1191],seed[3003],seed[873],seed[1384],seed[668],seed[91],seed[2724],seed[213],seed[136],seed[3179],seed[2537],seed[3588],seed[3306],seed[134],seed[3536],seed[4031],seed[3576],seed[4013],seed[4034],seed[2112],seed[3770],seed[2276],seed[1736],seed[1673],seed[2325],seed[2185],seed[334],seed[1389],seed[1853],seed[2865],seed[1168],seed[730],seed[1758],seed[930],seed[2347],seed[2096],seed[1445],seed[3436],seed[3061],seed[3119],seed[3029],seed[1761],seed[1824],seed[3191],seed[2099],seed[2882],seed[3554],seed[1010],seed[1422],seed[3847],seed[2673],seed[145],seed[1037],seed[814],seed[3447],seed[418],seed[2362],seed[1814],seed[1986],seed[2488],seed[2544],seed[2555],seed[3161],seed[695],seed[3803],seed[3513],seed[743],seed[57],seed[3096],seed[1122],seed[113],seed[879],seed[666],seed[1343],seed[3103],seed[3683],seed[2523],seed[400],seed[2706],seed[3756],seed[198],seed[1868],seed[594],seed[3299],seed[3485],seed[514],seed[3692],seed[1295],seed[1165],seed[571],seed[318],seed[2766],seed[716],seed[3723],seed[1113],seed[3944],seed[2711],seed[3437],seed[1753],seed[3917],seed[4030],seed[3377],seed[1320],seed[3304],seed[2501],seed[765],seed[1907],seed[464],seed[2468],seed[2159],seed[2162],seed[3972],seed[3663],seed[3137],seed[1234],seed[3604],seed[1912],seed[724],seed[1282],seed[4010],seed[1364],seed[806],seed[2180],seed[2177],seed[2691],seed[1794],seed[482],seed[3263],seed[43],seed[1609],seed[1110],seed[2271],seed[660],seed[2540],seed[164],seed[3149],seed[2876],seed[4038],seed[2749],seed[2443],seed[3186],seed[1917],seed[1226],seed[1303],seed[1382],seed[4083],seed[3247],seed[3725],seed[1978],seed[3799],seed[1663],seed[1963],seed[1661],seed[1173],seed[3389],seed[1084],seed[2379],seed[1548],seed[1581],seed[2140],seed[86],seed[2139],seed[1631],seed[1565],seed[1016],seed[3857],seed[1662],seed[669],seed[2593],seed[2235],seed[493],seed[1556],seed[3643],seed[1827],seed[203],seed[2971],seed[1882],seed[2573],seed[2729],seed[3388],seed[1008],seed[1820],seed[2105],seed[1604],seed[2286],seed[469],seed[2182],seed[1481],seed[1498],seed[3714],seed[1120],seed[2681],seed[821],seed[2457],seed[2369],seed[2830],seed[2841],seed[192],seed[3949],seed[2380],seed[3654],seed[2152],seed[788],seed[62],seed[424],seed[1945],seed[3537],seed[2174],seed[121],seed[1731],seed[1769],seed[2024],seed[4028],seed[779],seed[3500],seed[3095],seed[1338],seed[2792],seed[3568],seed[2220],seed[294],seed[3259],seed[3580],seed[2966],seed[3469],seed[2224],seed[593],seed[2259],seed[163],seed[4029],seed[89],seed[635],seed[2814],seed[1648],seed[3664],seed[1686],seed[501],seed[2028],seed[2644],seed[3367],seed[398],seed[179],seed[4036],seed[2114],seed[2700],seed[1681],seed[2211],seed[1124],seed[218],seed[961],seed[1603],seed[1576],seed[4033],seed[32],seed[1810],seed[710],seed[1523],seed[3081],seed[2538],seed[3769],seed[1036],seed[2254],seed[331],seed[619],seed[1747],seed[1231],seed[916],seed[2810],seed[670],seed[2856],seed[2909],seed[2989],seed[3833],seed[1552],seed[1875],seed[3657],seed[153],seed[1887],seed[2845],seed[2189],seed[2396],seed[119],seed[1247],seed[2258],seed[1239],seed[897],seed[1167],seed[27],seed[2352],seed[1732],seed[1668],seed[4079],seed[866],seed[376],seed[280],seed[3570],seed[224],seed[2109],seed[64],seed[2634],seed[764],seed[1733],seed[401],seed[3392],seed[2799],seed[2252],seed[3370],seed[1694],seed[663],seed[2102],seed[3650],seed[1171],seed[715],seed[2355],seed[4000],seed[1403],seed[1327],seed[2419],seed[1192],seed[3176],seed[3118],seed[4061],seed[667],seed[2956],seed[1594],seed[292],seed[3348],seed[2010],seed[2866],seed[2979],seed[2015],seed[3625],seed[3285],seed[3087],seed[2715],seed[3281],seed[546],seed[974],seed[1372],seed[438],seed[82],seed[3257],seed[1209],seed[1608],seed[1563],seed[3746],seed[758],seed[991],seed[40],seed[1539],seed[2798],seed[259],seed[1223],seed[2770],seed[3704],seed[3516],seed[1236],seed[2855],seed[2366],seed[3503],seed[3380],seed[2322],seed[1190],seed[78],seed[3262],seed[2414],seed[2565],seed[295],seed[2977],seed[2237],seed[527],seed[3786],seed[605],seed[2887],seed[1118],seed[3312],seed[1104],seed[2788],seed[1995],seed[3738],seed[3473],seed[494],seed[1803],seed[440],seed[1513],seed[746],seed[628],seed[177],seed[1428],seed[1509],seed[1194],seed[2201],seed[329],seed[2209],seed[574],seed[2067],seed[3470],seed[3563],seed[4068],seed[834],seed[3703],seed[775],seed[485],seed[1324],seed[322],seed[3239],seed[836],seed[3638],seed[30],seed[303],seed[45],seed[2852],seed[542],seed[944],seed[1629],seed[721],seed[2327],seed[2062],seed[1611],seed[2359],seed[1479],seed[3241],seed[862],seed[3812],seed[1956],seed[649],seed[793],seed[596],seed[2508],seed[1164],seed[3078],seed[2778],seed[899],seed[3159],seed[3674],seed[1186],seed[2312],seed[1800],seed[1780],seed[1806],seed[478],seed[1813],seed[142],seed[2692],seed[1898],seed[371],seed[3932],seed[2372],seed[3424],seed[1248],seed[2090],seed[31],seed[1957],seed[3223],seed[2316],seed[1116],seed[2833],seed[4059],seed[1616],seed[1289],seed[2331],seed[3073],seed[3816],seed[1701],seed[1526],seed[508],seed[1462],seed[2986],seed[3493],seed[2763],seed[2846],seed[3108],seed[3060],seed[364],seed[982],seed[2350],seed[3656],seed[2987],seed[3755],seed[1591],seed[1979],seed[2313],seed[1106],seed[2748],seed[1589],seed[599],seed[2421],seed[3566],seed[3871],seed[3353],seed[1408],seed[932],seed[3475],seed[2405],seed[3144],seed[3162],seed[439],seed[308],seed[2955],seed[3154],seed[2704],seed[23],seed[3877],seed[3922],seed[2019],seed[1825],seed[72],seed[1799],seed[1586],seed[1497],seed[893],seed[2040],seed[36],seed[16],seed[1053],seed[3236],seed[2886],seed[654],seed[519],seed[2155],seed[2607],seed[346],seed[818],seed[1334],seed[39],seed[831],seed[407],seed[1101],seed[1238],seed[309],seed[1697],seed[1281],seed[3868],seed[1561],seed[3422],seed[2226],seed[1724],seed[3310],seed[855],seed[622],seed[3763],seed[3194],seed[3822],seed[1176],seed[2740],seed[433],seed[3810],seed[2144],seed[518],seed[1227],seed[3052],seed[2374],seed[3411],seed[109],seed[1260],seed[284],seed[1347],seed[3220],seed[392],seed[3440],seed[1169],seed[1270],seed[1626],seed[1968],seed[645],seed[3244],seed[2579],seed[2032],seed[1336],seed[911],seed[2427],seed[1850],seed[3334],seed[2602],seed[1804],seed[1764],seed[2239],seed[979],seed[2975],seed[2650],seed[2600],seed[2877],seed[1961],seed[2231],seed[2831],seed[2121],seed[1012],seed[41],seed[233],seed[2341],seed[3338],seed[3288],seed[1551],seed[1880],seed[3775],seed[2589],seed[1743],seed[3669],seed[1383],seed[1905],seed[3827],seed[537],seed[2036],seed[3442],seed[310],seed[2458],seed[281],seed[2658],seed[1700],seed[3023],seed[3887],seed[884],seed[3099],seed[3115],seed[3234],seed[361],seed[399],seed[3013],seed[3265],seed[1319],seed[2726],seed[3726],seed[2416],seed[1357],seed[1066],seed[2980],seed[208],seed[1580],seed[3771],seed[3975],seed[52],seed[154],seed[3342],seed[2305],seed[3564],seed[2007],seed[1935],seed[547],seed[3924],seed[2335],seed[769],seed[1096],seed[3992],seed[1391],seed[920],seed[2320],seed[2969],seed[1043],seed[1099],seed[2490],seed[2874],seed[2170],seed[2598],seed[3521],seed[3021],seed[1271],seed[3336],seed[4053],seed[1989],seed[3860],seed[2],seed[590],seed[3599],seed[2561],seed[1822],seed[2758],seed[2065],seed[1547],seed[3603],seed[252],seed[3789],seed[1444],seed[1107],seed[1291],seed[1442],seed[2329],seed[456],seed[2398],seed[2401],seed[3344],seed[2623],seed[540],seed[2652],seed[3136],seed[1143],seed[3911],seed[1953],seed[3546],seed[1405],seed[38],seed[3686],seed[3595],seed[3350],seed[1103],seed[2008],seed[1578],seed[1419],seed[20],seed[3920],seed[2656],seed[3100],seed[1177],seed[2664],seed[3814],seed[3904],seed[155],seed[3742],seed[1235],seed[4069],seed[170],seed[2851],seed[3421],seed[390],seed[2097],seed[3477],seed[1900],seed[2686],seed[3508],seed[1006],seed[3123],seed[4023],seed[2592],seed[772],seed[3152],seed[3291],seed[277],seed[3862],seed[3826],seed[235],seed[3056],seed[1432],seed[263],seed[852],seed[3232],seed[871],seed[239],seed[3148],seed[1997],seed[2038],seed[262],seed[2358],seed[790],seed[1531],seed[832],seed[967],seed[161],seed[93],seed[858],seed[111],seed[840],seed[475],seed[985],seed[2645],seed[1973],seed[2225],seed[3700],seed[3606],seed[2440],seed[144],seed[2265],seed[3600],seed[3107],seed[3733],seed[3720],seed[3907],seed[3360],seed[3098],seed[483],seed[1454],seed[2564],seed[881],seed[4052],seed[621],seed[506],seed[800],seed[2476],seed[3804],seed[3160],seed[921],seed[1204],seed[889],seed[1575],seed[1083],seed[910],seed[2871],seed[3979],seed[701],seed[2993],seed[1750],seed[2382],seed[2207],seed[1839],seed[221],seed[1172],seed[3569],seed[1155],seed[42],seed[2803],seed[498],seed[1632],seed[3721],seed[1902],seed[3460],seed[50],seed[2275],seed[2486],seed[2849],seed[386],seed[397],seed[338],seed[2878],seed[2368],seed[234],seed[2394],seed[1467],seed[1914],seed[822],seed[2637],seed[54],seed[195],seed[1095],seed[5],seed[1706],seed[1022],seed[2697],seed[3126],seed[3416],seed[3201],seed[2281],seed[1128],seed[4041],seed[2868],seed[3138],seed[12],seed[1828],seed[1407],seed[2937],seed[1994],seed[983],seed[528],seed[2266],seed[2694],seed[1675],seed[3954],seed[1719],seed[2586],seed[2869],seed[2083],seed[1390],seed[1693],seed[3623],seed[2387],seed[2822],seed[2791],seed[3925],seed[3559],seed[3233],seed[2111],seed[630],seed[2365],seed[581],seed[1480],seed[3929],seed[1550],seed[1981],seed[1582],seed[3200],seed[2893],seed[739],seed[3212],seed[3357],seed[1643],seed[3910],seed[3133],seed[1314],seed[3207],seed[895],seed[2604],seed[2647],seed[3520],seed[3523],seed[1417],seed[2982],seed[802],seed[850],seed[1845],seed[3943],seed[2924],seed[2053],seed[2479],seed[2773],seed[939],seed[3959],seed[3020],seed[3203],seed[3278],seed[532],seed[2743],seed[2296],seed[653],seed[3110],seed[1704],seed[2370],seed[349],seed[2236],seed[266],seed[1698],seed[567],seed[2742],seed[3737],seed[3611],seed[3633],seed[2525],seed[507],seed[3174],seed[3675],seed[129],seed[3292],seed[990],seed[2444],seed[1274],seed[2092],seed[2198],seed[317],seed[914],seed[3927],seed[3289],seed[1938],seed[2156],seed[2208],seed[3648],seed[2663],seed[118],seed[4060],seed[1932],seed[2927],seed[942],seed[1773],seed[3318],seed[887],seed[1528],seed[545],seed[2826],seed[196],seed[3129],seed[1212],seed[2705],seed[2137],seed[1061],seed[2885],seed[2353],seed[2172],seed[1218],seed[791],seed[1862],seed[1711],seed[207],seed[3498],seed[3075],seed[4076],seed[1566],seed[3937],seed[784],seed[1351],seed[2079],seed[1713],seed[1206],seed[3875],seed[412],seed[3373],seed[2255],seed[2653],seed[3219],seed[1888],seed[577],seed[3684],seed[1368],seed[2035],seed[4082],seed[2084],seed[1406],seed[3143],seed[3048],seed[3915],seed[3482],seed[3958],seed[4075],seed[2786],seed[3158],seed[2670],seed[3779],seed[1756],seed[232],seed[601],seed[3337],seed[1263],seed[2765],seed[924],seed[1353],seed[711],seed[3728],seed[2157],seed[34],seed[2323],seed[44],seed[568],seed[3572],seed[2923],seed[51],seed[2491],seed[1471],seed[2717],seed[447],seed[708],seed[2668],seed[1046],seed[2200],seed[820],seed[1105],seed[1376],seed[2059],seed[3466],seed[1504],seed[2601],seed[2044],seed[3586],seed[1919],seed[808],seed[3109],seed[2796],seed[3928],seed[3767],seed[4080],seed[2737],seed[100],seed[2671],seed[1415],seed[2408],seed[3311],seed[1094],seed[1305],seed[2230],seed[1505],seed[2435],seed[465],seed[3781],seed[4009],seed[4086],seed[778],seed[2418],seed[640],seed[2500],seed[2025],seed[257],seed[2662],seed[2720],seed[267],seed[2582],seed[625],seed[2958],seed[3055],seed[2166],seed[3912],seed[1033],seed[3049],seed[2847],seed[3501],seed[1714],seed[3349],seed[1771],seed[3828],seed[1076],seed[3333],seed[3268],seed[584],seed[1004],seed[468],seed[1111],seed[2646],seed[1625],seed[2591],seed[682],seed[2424],seed[1117],seed[1495],seed[497],seed[890],seed[993],seed[2547],seed[610],seed[526],seed[472],seed[328],seed[865],seed[3544],seed[11],seed[3214],seed[2354],seed[3825],seed[87],seed[1795],seed[3031],seed[432],seed[2782],seed[1035],seed[1379],seed[1257],seed[21],seed[3558],seed[2665],seed[3346],seed[647],seed[1203],seed[946],seed[3015],seed[1125],seed[2516],seed[3791],seed[1411],seed[2227],seed[2006],seed[2921],seed[1399],seed[984],seed[3017],seed[3978],seed[3301],seed[2639],seed[3208],seed[220],seed[935],seed[3705],seed[1311],seed[3639],seed[3869],seed[2640],seed[566],seed[1687],seed[755],seed[365],seed[1569],seed[1722],seed[2840],seed[2961],seed[740],seed[559],seed[1214],seed[3374],seed[2914],seed[3303],seed[579],seed[796],seed[4004],seed[2524],seed[3973],seed[353],seed[479],seed[1876],seed[3340],seed[1646],seed[3205],seed[2428],seed[1808],seed[413],seed[612],seed[1443],seed[1606],seed[1744],seed[573],seed[3282],seed[2480],seed[2781],seed[1717],seed[1396],seed[3524],seed[332],seed[101],seed[3735],seed[713],seed[2575],seed[1983],seed[1819],seed[1929],seed[3963],seed[2628],seed[664],seed[2103],seed[725],seed[313],seed[1222],seed[2896],seed[3512],seed[1063],seed[3326],seed[2195],seed[2735],seed[1229],seed[2318],seed[2535],seed[4019],seed[421],seed[3171],seed[587],seed[2232],seed[4040],seed[249],seed[2635],seed[58],seed[3903],seed[2970],seed[306],seed[2357],seed[3853],seed[1931],seed[2453],seed[2193],seed[405],seed[1924],seed[3831],seed[637],seed[2873],seed[3204],seed[2513],seed[1520],seed[2000],seed[1494],seed[2509],seed[219],seed[2505],seed[3731],seed[1491],seed[3696],seed[1921],seed[94],seed[3790],seed[359],seed[4064],seed[356],seed[2917],seed[448],seed[1967],seed[2619],seed[2315],seed[2819],seed[1805],seed[449],seed[1508],seed[908],seed[3764],seed[1097],seed[1300],seed[512],seed[958],seed[1934],seed[360],seed[2689],seed[2913],seed[4074],seed[810],seed[2441],seed[1482],seed[1834],seed[774],seed[2406],seed[73],seed[894],seed[1323],seed[2074],seed[1423],seed[2801],seed[4039],seed[804],seed[97],seed[417],seed[575],seed[1776],seed[2562],seed[3793],seed[2397],seed[1607],seed[3252],seed[1426],seed[2095],seed[2859],seed[2702],seed[3849],seed[59],seed[2214],seed[3238],seed[1889],seed[3381],seed[617],seed[228],seed[1048],seed[904],seed[1702],seed[2392],seed[2787],seed[2395],seed[7],seed[2284],seed[3981],seed[1065],seed[1202],seed[261],seed[1242],seed[2212],seed[1028],seed[3140],seed[1506],seed[15],seed[131],seed[2587],seed[3716],seed[3815],seed[1210],seed[287],seed[520],seed[1127],seed[395],seed[2596],seed[1980],seed[684],seed[2243],seed[1185],seed[704],seed[2233],seed[2930],seed[2655],seed[1510],seed[1250],seed[3276],seed[1703],seed[1093],seed[1340],seed[3113],seed[1425],seed[905],seed[251],seed[2013],seed[797],seed[4062],seed[675],seed[3708],seed[3717],seed[1418],seed[2660],seed[2529],seed[3998],seed[1843],seed[3022],seed[1883],seed[3286],seed[3451],seed[4015],seed[3578],seed[2364],seed[2273],seed[2947],seed[3834],seed[1148],seed[2627],seed[3551],seed[3821],seed[1707],seed[3990],seed[642],seed[1901],seed[137],seed[46],seed[1585],seed[1],seed[138],seed[1972],seed[2106],seed[2247],seed[1705],seed[1587],seed[3322],seed[1903],seed[2039],seed[687],seed[451],seed[2135],seed[1628],seed[2848],seed[3867],seed[1998],seed[3327],seed[2542],seed[2082],seed[3722],seed[2978],seed[2614],seed[2824],seed[236],seed[1346],seed[484],seed[1108],seed[934],seed[1507],seed[877],seed[3997],seed[2780],seed[1013],seed[1775],seed[3405],seed[583],seed[2557],seed[2223],seed[901],seed[3807],seed[2113],seed[2836],seed[3976],seed[1365],seed[3266],seed[947],seed[3053],seed[922],seed[4037],seed[3293],seed[1249],seed[0],seed[2821],seed[354],seed[1069],seed[70],seed[3908],seed[2922],seed[1071],seed[76],seed[1777],seed[2863],seed[2757],seed[1672],seed[3898],seed[773],seed[2014],seed[888],seed[3951],seed[2680],seed[480],seed[1562],seed[2775],seed[2620],seed[3690],seed[1306],seed[2433],seed[3715],seed[1301],seed[3251],seed[677],seed[3739],seed[691],seed[2825],seed[319],seed[3662],seed[1666],seed[1598],seed[3581],seed[245],seed[2744],seed[2963],seed[314],seed[727],seed[387],seed[3845],seed[3858],seed[124],seed[4048],seed[3316],seed[4092],seed[114],seed[1394],seed[1676],seed[948],seed[604],seed[2104],seed[678],seed[1219],seed[68],seed[2910],seed[436],seed[2404],seed[3514],seed[3574],seed[1044],seed[1355],seed[2533],seed[1635],seed[1765],seed[2651],seed[3216],seed[3481],seed[133],seed[2291],seed[3454],seed[925],seed[339],seed[2009],seed[3748],seed[3438],seed[3863],seed[3283],seed[3605],seed[3744],seed[4066],seed[2016],seed[2528],seed[1590],seed[2998],seed[430],seed[733],seed[1246],seed[2438],seed[466],seed[286],seed[950],seed[513],seed[3632],seed[544],seed[3953],seed[2240],seed[2768],seed[1068],seed[2837],seed[1788],seed[3582],seed[1533],seed[2738],seed[3819],seed[1554],seed[2552],seed[700],seed[3471],seed[2384],seed[2531],seed[156],seed[3947],seed[2512],seed[422],seed[3260],seed[1266],seed[1944],seed[1653],seed[3499],seed[3601],seed[3444],seed[2021],seed[272],seed[3977],seed[4024],seed[2806],seed[1361],seed[4047],seed[2594],seed[3321],seed[3014],seed[2566],seed[1280],seed[2439],seed[3284],seed[2116],seed[3938],seed[3967],seed[1472],seed[569],seed[1091],seed[3125],seed[250],seed[3489],seed[325],seed[2940],seed[1774],seed[633],seed[815],seed[657],seed[1080],seed[3565],seed[1252],seed[3874],seed[2649],seed[2879],seed[2378],seed[1996],seed[2809],seed[1784],seed[2376],seed[385],seed[745],seed[1659],seed[3542],seed[2942],seed[388],seed[2334],seed[1863],seed[2075],seed[3305],seed[199],seed[3956],seed[3324],seed[3426],seed[1618],seed[636],seed[2741],seed[3192],seed[2794],seed[2807],seed[3261],seed[211],seed[3449],seed[2590],seed[226],seed[2974],seed[4027],seed[1436],seed[688],seed[1187],seed[2093],seed[886],seed[2017],seed[638],seed[1160],seed[1448],seed[3480],seed[3842],seed[2759],seed[3617],seed[505],seed[3227],seed[980],seed[3724],seed[1920],seed[183],seed[2559],seed[1891],seed[414],seed[3045],seed[1197],seed[215],seed[523],seed[3987],seed[1864],seed[702],seed[2115],seed[3671],seed[3890],seed[1682],seed[3864],seed[854],seed[3758],seed[3999],seed[348],seed[1660],seed[2260],seed[3667],seed[3106],seed[641],seed[1182],seed[9],seed[1851],seed[3390],seed[3196],seed[994],seed[1742],seed[2659],seed[151],seed[446],seed[1163],seed[3250],seed[3850],seed[845],seed[1149],seed[99],seed[3494],seed[535],seed[4055],seed[1142],seed[876],seed[2904],seed[2581],seed[2756],seed[728],seed[3141],seed[1692],seed[143],seed[1283],seed[798],seed[1030],seed[825],seed[1958],seed[3994],seed[2420],seed[10],seed[2011],seed[3150],seed[3050],seed[1304],seed[3934],seed[941],seed[186],seed[463],seed[1050],seed[1134],seed[3294],seed[870],seed[394],seed[3047],seed[1881],seed[3697],seed[3772],seed[24],seed[3461],seed[3147],seed[578],seed[735],seed[3743],seed[268],seed[1179],seed[753],seed[2409],seed[1842],seed[2818],seed[2920],seed[1915],seed[3044],seed[951],seed[2599],seed[2550],seed[1077],seed[2746],seed[3950],seed[3464],seed[2188],seed[3298],seed[3005],seed[355],seed[2244],seed[320],seed[2125],seed[3507],seed[3622],seed[2603],seed[1529],seed[290],seed[1031],seed[389],seed[1751],seed[2745],seed[3386],seed[3274],seed[1089],seed[1966],seed[616],seed[1354],seed[1976],seed[492],seed[1253],seed[1489],seed[160],seed[1318],seed[792],seed[1927],seed[2326],seed[2929],seed[147],seed[1477],seed[162],seed[2954],seed[2173],seed[2375],seed[1385],seed[757],seed[923],seed[3018],seed[699],seed[1100],seed[382],seed[3627],seed[3],seed[141],seed[3980],seed[2431],seed[293],seed[248],seed[1540],seed[3366],seed[3996],seed[1783],seed[2460],seed[3335],seed[883],seed[843],seed[1441],seed[842],seed[25],seed[3414],seed[3844],seed[1375],seed[4006],seed[2817],seed[977],seed[867],seed[122],seed[1402],seed[2951],seed[1456],seed[1470],seed[1519],seed[3515],seed[2892],seed[79],seed[3183],seed[1287],seed[1421],seed[1787],seed[3762],seed[2793],seed[3146],seed[1137],seed[3813],seed[2721],seed[3691],seed[525],seed[789],seed[1535],seed[998],seed[1193],seed[1930],seed[2518],seed[247],seed[1367],seed[844],seed[1156],seed[1259],seed[1434],seed[2907],seed[214],seed[2795],seed[1207],seed[3290],seed[1486],seed[1189],seed[375],seed[2089],seed[1377],seed[819],seed[2131],seed[2567],seed[315],seed[3228],seed[3945],seed[3030],seed[3368],seed[1559],seed[3072],seed[3802],seed[970],seed[3213],seed[2727],seed[2150],seed[1151],seed[2217],seed[2761],seed[2306],seed[3619],seed[3525],seed[812],seed[2965],seed[3809],seed[754],seed[709],seed[1789],seed[2194],seed[3432],seed[2151],seed[4018],seed[2953],seed[270],seed[458],seed[1397],seed[1251],seed[3694],seed[3175],seed[1288],seed[2219],seed[3242],seed[1597],seed[2883],seed[1835],seed[3902],seed[1041],seed[159],seed[1564],seed[1951],seed[460],seed[2832],seed[229],seed[1993],seed[3651],seed[3474],seed[81],seed[3124],seed[2931],seed[3385],seed[202],seed[3193],seed[2530],seed[330],seed[3173],seed[3038],seed[777],seed[959],seed[2060],seed[3545],seed[3916],seed[3888],seed[2447],seed[2342],seed[2402],seed[694],seed[2919],seed[1943],seed[1115],seed[2383],seed[1290],seed[1797],seed[3006],seed[3666],seed[2410],seed[321],seed[8],seed[4078],seed[1284],seed[3468],seed[2091],seed[3296],seed[1315],seed[1849],seed[1329],seed[2585],seed[1199],seed[3532],seed[2597],seed[2895],seed[2783],seed[1837],seed[976],seed[2981],seed[693],seed[84],seed[1815],seed[1216],seed[2241],seed[3594],seed[966],seed[2685],seed[1757],seed[3084],seed[554],seed[3843],seed[661],seed[370],seed[1332],seed[4012],seed[307],seed[1232],seed[3805],seed[2330],seed[3398],seed[3538],seed[489],seed[2834],seed[591],seed[1420],seed[1522],seed[3923],seed[570],seed[3248],seed[551],seed[470],seed[2541],seed[416],seed[2912],seed[1844],seed[3448],seed[2677],seed[326],seed[3164],seed[1485],seed[2842],seed[1859],seed[2838],seed[102],seed[3307],seed[3540],seed[937],seed[3754],seed[3382],seed[2606],seed[2204],seed[720],seed[1946],seed[4007],seed[2087],seed[2210],seed[2771],seed[3837],seed[1671],seed[783],seed[1090],seed[408],seed[3612],seed[2388],seed[3425],seed[2933],seed[1879],seed[3051],seed[2202],seed[2894],seed[2169],seed[2454],seed[3901],seed[3679],seed[2915],seed[690],seed[3882],seed[1553],seed[3955],seed[3552],seed[74],seed[3273],seed[1058],seed[1447],seed[172],seed[1401],seed[2412],seed[1009],seed[809],seed[3510],seed[2455],seed[3046],seed[3982],seed[3750],seed[3231],seed[2456],seed[2959],seed[872],seed[3415],seed[140],seed[1294],seed[1892],seed[2287],seed[175],seed[3035],seed[1909],seed[3184],seed[3644],seed[1224],seed[3401],seed[296],seed[369],seed[762],seed[683],seed[312],seed[1541],seed[3593],seed[3443],seed[3689],seed[1992],seed[1060],seed[564],seed[3456],seed[1624],seed[536],seed[3590],seed[1877],seed[278],seed[3765],seed[3682],seed[1831],seed[2957],seed[2348],seed[2493],seed[3711],seed[1166],seed[2127],seed[3300],seed[1767],seed[1527]}),
        .cross_prob(cross_prob),
        .codeword(codeword8),
        .received(received8)
        );
    
    bsc bsc9(
        .clk(clk),
        .reset(reset),
        .seed({seed[260],seed[737],seed[3850],seed[3852],seed[2184],seed[422],seed[1938],seed[626],seed[753],seed[3877],seed[522],seed[4011],seed[60],seed[3657],seed[1669],seed[2945],seed[549],seed[1798],seed[3738],seed[2443],seed[2663],seed[2384],seed[851],seed[2015],seed[1088],seed[2265],seed[472],seed[1429],seed[1388],seed[2101],seed[3797],seed[3687],seed[946],seed[1090],seed[3151],seed[749],seed[262],seed[464],seed[747],seed[294],seed[3960],seed[672],seed[2219],seed[3893],seed[1908],seed[3924],seed[3750],seed[1568],seed[67],seed[3965],seed[3925],seed[1361],seed[536],seed[4084],seed[3574],seed[2701],seed[17],seed[820],seed[3895],seed[78],seed[2657],seed[2516],seed[321],seed[2159],seed[284],seed[392],seed[568],seed[2831],seed[1614],seed[2951],seed[1706],seed[3890],seed[1073],seed[1877],seed[1322],seed[771],seed[1256],seed[3918],seed[1271],seed[3961],seed[1081],seed[3222],seed[3365],seed[1895],seed[2475],seed[1520],seed[1664],seed[3744],seed[3701],seed[3772],seed[2827],seed[145],seed[1534],seed[223],seed[920],seed[3449],seed[4043],seed[1215],seed[2463],seed[3028],seed[2422],seed[230],seed[2494],seed[10],seed[1760],seed[2865],seed[2111],seed[1393],seed[1161],seed[3620],seed[3366],seed[871],seed[2260],seed[1855],seed[2414],seed[19],seed[4069],seed[3352],seed[1213],seed[1439],seed[1503],seed[163],seed[1363],seed[3896],seed[3052],seed[2278],seed[693],seed[1681],seed[526],seed[1595],seed[240],seed[809],seed[2526],seed[383],seed[2741],seed[1484],seed[2661],seed[2224],seed[80],seed[151],seed[1633],seed[2832],seed[1644],seed[1368],seed[832],seed[1165],seed[3327],seed[277],seed[3729],seed[1238],seed[416],seed[181],seed[1015],seed[2479],seed[106],seed[573],seed[3667],seed[810],seed[1834],seed[252],seed[1533],seed[2651],seed[3886],seed[484],seed[2131],seed[2783],seed[3487],seed[927],seed[1913],seed[1299],seed[2193],seed[382],seed[577],seed[118],seed[160],seed[1536],seed[2570],seed[2162],seed[479],seed[2069],seed[2989],seed[990],seed[1601],seed[3663],seed[1784],seed[2816],seed[2204],seed[3868],seed[2615],seed[885],seed[33],seed[2133],seed[2825],seed[3074],seed[1233],seed[1797],seed[1637],seed[4028],seed[2],seed[1435],seed[2129],seed[2499],seed[1096],seed[1738],seed[4068],seed[2503],seed[2396],seed[1675],seed[3742],seed[2483],seed[2359],seed[1773],seed[958],seed[3548],seed[1485],seed[1505],seed[1867],seed[3575],seed[2685],seed[1692],seed[3088],seed[9],seed[1655],seed[3811],seed[3810],seed[410],seed[2586],seed[1795],seed[3677],seed[2058],seed[1274],seed[760],seed[2904],seed[3529],seed[1513],seed[3482],seed[1626],seed[3038],seed[4080],seed[451],seed[698],seed[1310],seed[2502],seed[3165],seed[3872],seed[2141],seed[1323],seed[1390],seed[4021],seed[3361],seed[485],seed[2279],seed[2137],seed[3375],seed[1830],seed[2621],seed[3532],seed[1980],seed[3188],seed[1995],seed[714],seed[2839],seed[1351],seed[2815],seed[1979],seed[3398],seed[3658],seed[650],seed[2342],seed[2769],seed[489],seed[649],seed[2188],seed[1755],seed[1904],seed[121],seed[3261],seed[278],seed[3536],seed[1244],seed[783],seed[2729],seed[3702],seed[2256],seed[1703],seed[1756],seed[3335],seed[4083],seed[2763],seed[2361],seed[584],seed[2940],seed[1540],seed[1531],seed[2715],seed[811],seed[4085],seed[1075],seed[114],seed[1879],seed[854],seed[470],seed[3178],seed[2071],seed[1967],seed[2233],seed[4042],seed[1432],seed[2863],seed[3565],seed[1635],seed[2976],seed[476],seed[1964],seed[3061],seed[3369],seed[2728],seed[3220],seed[1340],seed[3092],seed[458],seed[2937],seed[2164],seed[667],seed[1001],seed[2477],seed[2762],seed[3413],seed[1929],seed[2196],seed[3539],seed[1229],seed[241],seed[1246],seed[1091],seed[957],seed[2946],seed[2488],seed[1876],seed[3740],seed[558],seed[2998],seed[1652],seed[1744],seed[882],seed[2645],seed[1304],seed[3727],seed[963],seed[3237],seed[1791],seed[92],seed[828],seed[2883],seed[3623],seed[887],seed[168],seed[499],seed[2474],seed[3119],seed[784],seed[2625],seed[1032],seed[2294],seed[4001],seed[3819],seed[3731],seed[726],seed[895],seed[245],seed[3224],seed[2211],seed[1611],seed[1321],seed[3],seed[388],seed[3194],seed[888],seed[3116],seed[3477],seed[1324],seed[3820],seed[3919],seed[994],seed[1739],seed[561],seed[1440],seed[542],seed[3948],seed[447],seed[2126],seed[3517],seed[1976],seed[1653],seed[563],seed[1122],seed[2482],seed[3084],seed[2374],seed[3436],seed[2817],seed[1730],seed[2529],seed[3757],seed[775],seed[3673],seed[1114],seed[2630],seed[567],seed[1647],seed[3916],seed[578],seed[3018],seed[2023],seed[425],seed[3577],seed[2844],seed[983],seed[1905],seed[2811],seed[3030],seed[759],seed[135],seed[1222],seed[4076],seed[3378],seed[3244],seed[1826],seed[2280],seed[2272],seed[3370],seed[3755],seed[681],seed[3037],seed[1582],seed[4022],seed[1207],seed[1950],seed[1766],seed[265],seed[3021],seed[1326],seed[655],seed[1139],seed[1620],seed[3474],seed[3480],seed[1731],seed[81],seed[2067],seed[2173],seed[2986],seed[2717],seed[2978],seed[3356],seed[2424],seed[1214],seed[4059],seed[3869],seed[2183],seed[2814],seed[2033],seed[2400],seed[841],seed[3763],seed[593],seed[3121],seed[270],seed[376],seed[3478],seed[2758],seed[1954],seed[924],seed[2476],seed[1859],seed[632],seed[24],seed[1226],seed[2754],seed[3271],seed[778],seed[3345],seed[1060],seed[3063],seed[3388],seed[870],seed[1374],seed[2478],seed[481],seed[1005],seed[2045],seed[3215],seed[452],seed[580],seed[620],seed[1162],seed[1003],seed[1259],seed[1893],seed[3911],seed[3341],seed[1850],seed[3706],seed[1423],seed[1287],seed[1919],seed[2667],seed[1884],seed[487],seed[3156],seed[740],seed[3445],seed[950],seed[3697],seed[1133],seed[2764],seed[1537],seed[1377],seed[2251],seed[2590],seed[930],seed[224],seed[3883],seed[1442],seed[1510],seed[674],seed[2709],seed[131],seed[1421],seed[2795],seed[562],seed[116],seed[507],seed[1254],seed[1932],seed[3363],seed[2725],seed[3389],seed[271],seed[2209],seed[285],seed[2680],seed[3636],seed[3174],seed[915],seed[772],seed[2852],seed[3837],seed[1205],seed[2270],seed[1914],seed[3198],seed[2934],seed[3241],seed[1977],seed[2489],seed[2267],seed[1722],seed[2583],seed[2650],seed[3679],seed[2303],seed[409],seed[3009],seed[3938],seed[3983],seed[2792],seed[492],seed[1149],seed[3200],seed[880],seed[897],seed[3932],seed[2580],seed[192],seed[362],seed[3034],seed[3199],seed[685],seed[3320],seed[724],seed[516],seed[1169],seed[607],seed[1425],seed[3471],seed[2659],seed[528],seed[2592],seed[4017],seed[1529],seed[3635],seed[3434],seed[1935],seed[1610],seed[3279],seed[3692],seed[389],seed[1911],seed[2755],seed[3977],seed[2149],seed[359],seed[253],seed[2076],seed[1196],seed[1695],seed[3336],seed[3264],seed[2561],seed[1105],seed[365],seed[3381],seed[4003],seed[341],seed[2991],seed[2740],seed[2223],seed[2089],seed[4053],seed[633],seed[328],seed[4044],seed[1415],seed[1183],seed[4012],seed[3722],seed[2871],seed[3280],seed[1565],seed[3934],seed[4052],seed[1912],seed[3286],seed[1454],seed[872],seed[1067],seed[2027],seed[2331],seed[611],seed[1062],seed[1087],seed[2026],seed[2834],seed[2555],seed[3664],seed[3616],seed[1378],seed[2077],seed[4073],seed[1843],seed[1632],seed[3380],seed[2882],seed[3265],seed[22],seed[1118],seed[1084],seed[764],seed[3631],seed[1143],seed[1469],seed[3659],seed[483],seed[2299],seed[1098],seed[1940],seed[3991],seed[2176],seed[1380],seed[2711],seed[3825],seed[105],seed[53],seed[838],seed[1209],seed[2011],seed[1342],seed[2138],seed[3922],seed[701],seed[1902],seed[1822],seed[2386],seed[1519],seed[3282],seed[3826],seed[3069],seed[3491],seed[2912],seed[1412],seed[3989],seed[503],seed[4078],seed[2720],seed[2132],seed[1587],seed[2339],seed[1414],seed[1251],seed[4082],seed[74],seed[3622],seed[3344],seed[873],seed[3598],seed[2369],seed[2050],seed[1449],seed[2212],seed[2931],seed[1642],seed[361],seed[457],seed[559],seed[2652],seed[1951],seed[3836],seed[3728],seed[1553],seed[3384],seed[218],seed[2771],seed[2363],seed[3470],seed[934],seed[411],seed[1943],seed[66],seed[85],seed[3259],seed[214],seed[101],seed[937],seed[1694],seed[3155],seed[3683],seed[2908],seed[1017],seed[3439],seed[3466],seed[4095],seed[736],seed[68],seed[490],seed[2139],seed[817],seed[312],seed[1571],seed[3218],seed[2406],seed[1556],seed[1934],seed[2087],seed[3442],seed[1494],seed[1372],seed[2693],seed[2648],seed[1008],seed[469],seed[2810],seed[3301],seed[2738],seed[3605],seed[3060],seed[2356],seed[1986],seed[2742],seed[1753],seed[2565],seed[344],seed[2522],seed[515],seed[2439],seed[3796],seed[807],seed[3905],seed[547],seed[2197],seed[2947],seed[2656],seed[1466],seed[2544],seed[3578],seed[2746],seed[1327],seed[2647],seed[2140],seed[2335],seed[2194],seed[2906],seed[3898],seed[3689],seed[1687],seed[1508],seed[1801],seed[505],seed[3624],seed[2036],seed[2282],seed[225],seed[1389],seed[1376],seed[1044],seed[1124],seed[1957],seed[1963],seed[1218],seed[1410],seed[1750],seed[149],seed[1330],seed[985],seed[2042],seed[619],seed[3912],seed[1134],seed[3000],seed[876],seed[72],seed[1135],seed[2995],seed[3937],seed[1997],seed[207],seed[1890],seed[1799],seed[2411],seed[1489],seed[329],seed[3660],seed[808],seed[2927],seed[3504],seed[696],seed[1184],seed[320],seed[1949],seed[1666],seed[1294],seed[3351],seed[1848],seed[834],seed[3047],seed[3584],seed[2423],seed[4050],seed[2856],seed[1206],seed[2128],seed[585],seed[2124],seed[3800],seed[3231],seed[795],seed[0],seed[502],seed[41],seed[1590],seed[2495],seed[973],seed[903],seed[126],seed[2387],seed[3230],seed[1194],seed[1593],seed[3748],seed[2878],seed[2498],seed[1718],seed[3402],seed[315],seed[812],seed[3394],seed[4051],seed[3254],seed[2899],seed[1999],seed[1459],seed[1433],seed[2547],seed[3817],seed[2599],seed[2365],seed[2596],seed[2239],seed[3208],seed[940],seed[3372],seed[1420],seed[3387],seed[3343],seed[902],seed[2035],seed[1464],seed[2727],seed[1998],seed[2925],seed[3016],seed[1982],seed[1178],seed[2576],seed[3779],seed[1186],seed[162],seed[2404],seed[3159],seed[3787],seed[1258],seed[2749],seed[2004],seed[3682],seed[1273],seed[442],seed[263],seed[430],seed[2905],seed[38],seed[3226],seed[2066],seed[1960],seed[694],seed[304],seed[1092],seed[3094],seed[951],seed[164],seed[700],seed[1463],seed[1093],seed[1418],seed[2012],seed[797],seed[923],seed[1193],seed[124],seed[20],seed[1262],seed[2354],seed[3073],seed[1020],seed[3596],seed[460],seed[2812],seed[2295],seed[2266],seed[1314],seed[2782],seed[3562],seed[420],seed[949],seed[2388],seed[3495],seed[3176],seed[2473],seed[3552],seed[2014],seed[314],seed[1255],seed[50],seed[2525],seed[1039],seed[529],seed[2722],seed[3758],seed[1926],seed[3297],seed[2465],seed[2790],seed[3821],seed[944],seed[517],seed[1146],seed[2710],seed[28],seed[1277],seed[3431],seed[2122],seed[441],seed[496],seed[2447],seed[3671],seed[3506],seed[2115],seed[1455],seed[1563],seed[2962],seed[1732],seed[3432],seed[3236],seed[519],seed[2921],seed[1985],seed[2930],seed[3847],seed[1891],seed[2459],seed[1574],seed[831],seed[996],seed[3319],seed[1608],seed[991],seed[2653],seed[981],seed[2043],seed[3309],seed[65],seed[3643],seed[2440],seed[1869],seed[3695],seed[3376],seed[2744],seed[3300],seed[3724],seed[3416],seed[1191],seed[1394],seed[3503],seed[712],seed[1269],seed[3425],seed[732],seed[4062],seed[426],seed[2671],seed[2629],seed[1270],seed[776],seed[814],seed[1079],seed[380],seed[2148],seed[2293],seed[2060],seed[3050],seed[1371],seed[2349],seed[4007],seed[2835],seed[2696],seed[2730],seed[3593],seed[3112],seed[2208],seed[2428],seed[2745],seed[3214],seed[2538],seed[3851],seed[1083],seed[1103],seed[1646],seed[676],seed[2956],seed[1402],seed[3813],seed[3433],seed[3401],seed[2130],seed[3240],seed[326],seed[35],seed[2171],seed[247],seed[189],seed[3429],seed[761],seed[1144],seed[2608],seed[1683],seed[4008],seed[2996],seed[555],seed[2971],seed[2517],seed[2773],seed[2959],seed[1847],seed[3579],seed[569],seed[3168],seed[1106],seed[1981],seed[2142],seed[3427],seed[237],seed[1082],seed[2275],seed[1373],seed[287],seed[2928],seed[3520],seed[1030],seed[2747],seed[1930],seed[208],seed[3806],seed[1672],seed[1689],seed[3903],seed[456],seed[1279],seed[1578],seed[1525],seed[3184],seed[2994],seed[3505],seed[3793],seed[1897],seed[1045],seed[1707],seed[1266],seed[122],seed[3901],seed[2924],seed[514],seed[369],seed[3457],seed[3681],seed[2378],seed[3367],seed[378],seed[3305],seed[1915],seed[3085],seed[2564],seed[3325],seed[550],seed[1509],seed[2330],seed[3324],seed[1275],seed[2532],seed[1102],seed[2665],seed[2784],seed[2367],seed[3071],seed[2724],seed[777],seed[4029],seed[2381],seed[1535],seed[953],seed[1132],seed[2602],seed[3939],seed[2200],seed[1638],seed[3914],seed[533],seed[434],seed[3768],seed[2167],seed[3990],seed[165],seed[1645],seed[2352],seed[2676],seed[2658],seed[234],seed[448],seed[258],seed[482],seed[2467],seed[413],seed[4049],seed[2048],seed[3762],seed[2344],seed[2981],seed[2416],seed[538],seed[715],seed[2348],seed[3417],seed[2531],seed[418],seed[3274],seed[589],seed[3861],seed[919],seed[2007],seed[3639],seed[1413],seed[1878],seed[2207],seed[662],seed[790],seed[3488],seed[911],seed[1263],seed[1684],seed[3233],seed[2796],seed[3680],seed[830],seed[1313],seed[2103],seed[2472],seed[3959],seed[1334],seed[2914],seed[1865],seed[1702],seed[3022],seed[2803],seed[1034],seed[242],seed[523],seed[2787],seed[4031],seed[1022],seed[1549],seed[2273],seed[3068],seed[874],seed[2262],seed[1078],seed[274],seed[3776],seed[3672],seed[1853],seed[2876],seed[232],seed[2707],seed[3360],seed[1941],seed[2415],seed[1058],seed[2125],seed[2420],seed[466],seed[146],seed[1029],seed[2751],seed[4040],seed[1828],seed[1174],seed[231],seed[2074],seed[1367],seed[4088],seed[3118],seed[1260],seed[1253],seed[613],seed[167],seed[1583],seed[669],seed[1825],seed[3704],seed[2743],seed[348],seed[3117],seed[183],seed[2603],seed[1631],seed[1910],seed[2307],seed[2366],seed[1267],seed[564],seed[4064],seed[3149],seed[371],seed[2896],seed[2395],seed[2999],seed[1806],seed[900],seed[2019],seed[444],seed[1970],seed[2527],seed[3334],seed[1043],seed[2198],seed[3694],seed[1216],seed[3947],seed[959],seed[1038],seed[762],seed[2988],seed[914],seed[3531],seed[73],seed[4077],seed[1307],seed[404],seed[3705],seed[3641],seed[1150],seed[3933],seed[2316],seed[2637],seed[1182],seed[2355],seed[1567],seed[2497],seed[3970],seed[3586],seed[236],seed[1456],seed[18],seed[1539],seed[3485],seed[2689],seed[2886],seed[3354],seed[3803],seed[2536],seed[2567],seed[3167],seed[638],seed[1800],seed[3467],seed[3113],seed[2687],seed[243],seed[3051],seed[3785],seed[2587],seed[1268],seed[1585],seed[2861],seed[3550],seed[1780],seed[2780],seed[4041],seed[2943],seed[1625],seed[4018],seed[36],seed[3899],seed[2859],seed[3346],seed[660],seed[2890],seed[3981],seed[1049],seed[3538],seed[4026],seed[3955],seed[3210],seed[3675],seed[2068],seed[799],seed[631],seed[2425],seed[431],seed[1765],seed[2860],seed[352],seed[1126],seed[741],seed[2543],seed[1396],seed[259],seed[658],seed[2813],seed[1618],seed[939],seed[1284],seed[63],seed[2686],seed[1077],seed[1002],seed[2049],seed[3067],seed[3368],seed[3272],seed[3311],seed[3713],seed[657],seed[1303],seed[3891],seed[2345],seed[868],seed[2059],seed[2391],seed[4009],seed[2110],seed[859],seed[3994],seed[3189],seed[1874],seed[3373],seed[787],seed[26],seed[1325],seed[3147],seed[1070],seed[3907],seed[3175],seed[3897],seed[1235],seed[1109],seed[1308],seed[3024],seed[1793],seed[3307],seed[1431],seed[863],seed[1783],seed[467],seed[2073],seed[2199],seed[134],seed[2634],seed[1486],seed[257],seed[2086],seed[1880],seed[1151],seed[3090],seed[2146],seed[974],seed[2627],seed[318],seed[3268],seed[2259],seed[3420],seed[3612],seed[791],seed[372],seed[2287],seed[52],seed[1315],seed[268],seed[2136],seed[1072],seed[1110],seed[908],seed[2308],seed[1329],seed[3594],seed[551],seed[144],seed[2703],seed[3095],seed[3227],seed[1318],seed[3143],seed[1434],seed[1054],seed[384],seed[898],seed[1492],seed[3732],seed[3963],seed[196],seed[1770],seed[471],seed[1408],seed[1860],seed[2786],seed[1286],seed[989],seed[3878],seed[3479],seed[1427],seed[2471],seed[2794],seed[600],seed[4061],seed[1570],seed[2119],seed[3743],seed[358],seed[1175],seed[248],seed[2096],seed[2848],seed[3291],seed[2206],seed[1426],seed[1713],seed[1691],seed[3603],seed[2550],seed[1842],seed[3871],seed[3041],seed[748],seed[4055],seed[2433],seed[594],seed[338],seed[2846],seed[636],seed[2549],seed[1771],seed[2523],seed[2179],seed[982],seed[2983],seed[2533],seed[1643],seed[3756],seed[3589],seed[3805],seed[414],seed[3975],seed[1648],seed[1397],seed[1239],seed[3475],seed[1548],seed[796],seed[2247],seed[1024],seed[2407],seed[119],seed[869],seed[2152],seed[3618],seed[2654],seed[2419],seed[689],seed[350],seed[999],seed[3968],seed[2158],seed[2877],seed[1208],seed[3760],seed[3749],seed[2768],seed[3980],seed[3554],seed[120],seed[1749],seed[1742],seed[3169],seed[1591],seed[2977],seed[2177],seed[355],seed[2394],seed[3129],seed[2808],seed[3486],seed[3696],seed[1579],seed[310],seed[1615],seed[3303],seed[2217],seed[3321],seed[449],seed[55],seed[3674],seed[148],seed[2009],seed[2697],seed[2845],seed[2975],seed[552],seed[1248],seed[1497],seed[1010],seed[3223],seed[279],seed[3128],seed[3927],seed[1152],seed[2150],seed[1560],seed[804],seed[3234],seed[3141],seed[2838],seed[1708],seed[2733],seed[157],seed[1907],seed[2958],seed[1623],seed[3322],seed[1789],seed[3708],seed[143],seed[826],seed[1354],seed[336],seed[1526],seed[319],seed[579],seed[850],seed[586],seed[2837],seed[2123],seed[190],seed[107],seed[351],seed[692],seed[1909],seed[3500],seed[6],seed[1296],seed[2559],seed[1820],seed[1942],seed[1052],seed[3876],seed[2098],seed[2143],seed[702],seed[3207],seed[3191],seed[3537],seed[2781],seed[23],seed[1019],seed[2281],seed[2001],seed[1220],seed[610],seed[3881],seed[91],seed[1341],seed[2120],seed[3515],seed[1515],seed[1659],seed[2153],seed[1063],seed[408],seed[4074],seed[3163],seed[1451],seed[3654],seed[3438],seed[3913],seed[3317],seed[2057],seed[1745],seed[3304],seed[1305],seed[2551],seed[971],seed[3638],seed[4067],seed[3684],seed[2731],seed[1348],seed[1725],seed[381],seed[2163],seed[1901],seed[3630],seed[3142],seed[1225],seed[2577],seed[3410],seed[3786],seed[544],seed[1831],seed[291],seed[878],seed[3070],seed[1465],seed[2085],seed[2867],seed[893],seed[1071],seed[665],seed[1792],seed[3172],seed[1617],seed[2225],seed[3610],seed[2759],seed[2623],seed[815],seed[2135],seed[3106],seed[1918],seed[104],seed[391],seed[2521],seed[1719],seed[1232],seed[504],seed[301],seed[948],seed[2232],seed[3145],seed[3996],seed[2181],seed[1927],seed[54],seed[246],seed[3754],seed[3296],seed[2093],seed[4],seed[518],seed[3784],seed[2668],seed[3295],seed[2493],seed[1285],seed[1845],seed[3774],seed[3422],seed[1966],seed[412],seed[2800],seed[1379],seed[2100],seed[402],seed[3253],seed[84],seed[3807],seed[3828],seed[1856],seed[2620],seed[4013],seed[141],seed[2038],seed[3374],seed[2913],seed[1882],seed[848],seed[2636],seed[3493],seed[1490],seed[3017],seed[1699],seed[2319],seed[677],seed[3588],seed[40],seed[3077],seed[2155],seed[2968],seed[3235],seed[705],seed[3508],seed[2005],seed[32],seed[2409],seed[1569],seed[2675],seed[3035],seed[76],seed[1155],seed[2664],seed[1572],seed[3428],seed[1336],seed[4015],seed[1829],seed[1530],seed[2606],seed[1042],seed[2041],seed[857],seed[2540],seed[3739],seed[3855],seed[896],seed[3252],seed[1355],seed[3582],seed[3686],seed[3213],seed[1074],seed[3138],seed[3476],seed[306],seed[2748],seed[309],seed[856],seed[2470],seed[781],seed[3250],seed[2210],seed[535],seed[3962],seed[1064],seed[2823],seed[2323],seed[446],seed[1844],seed[1243],seed[3652],seed[424],seed[1197],seed[1219],seed[3314],seed[2907],seed[531],seed[3201],seed[3444],seed[5],seed[169],seed[864],seed[3964],seed[3440],seed[3809],seed[2053],seed[2075],seed[2218],seed[918],seed[1991],seed[1817],seed[2866],seed[618],seed[1704],seed[1762],seed[2328],seed[4046],seed[1900],seed[3115],seed[1369],seed[763],seed[1236],seed[191],seed[3693],seed[2157],seed[98],seed[2973],seed[1366],seed[2916],seed[102],seed[295],seed[3802],seed[745],seed[3556],seed[2376],seed[1627],seed[2236],seed[2434],seed[174],seed[2510],seed[588],seed[933],seed[3735],seed[1339],seed[998],seed[548],seed[1931],seed[909],seed[1483],seed[798],seed[1224],seed[1240],seed[2254],seed[2405],seed[2195],seed[2901],seed[1794],seed[4072],seed[601],seed[2557],seed[1894],seed[226],seed[1381],seed[1417],seed[1297],seed[2088],seed[1682],seed[1737],seed[616],seed[1936],seed[390],seed[2604],seed[1823],seed[2230],seed[2134],seed[3928],seed[3759],seed[1883],seed[1457],seed[2456],seed[3604],seed[4086],seed[2888],seed[3353],seed[3882],seed[906],seed[3986],seed[3269],seed[1338],seed[3059],seed[1796],seed[766],seed[2505],seed[438],seed[3211],seed[1317],seed[1405],seed[3124],seed[3248],seed[2949],seed[500],seed[2034],seed[3019],seed[1157],seed[3350],seed[1899],seed[363],seed[2340],seed[2723],seed[3012],seed[3767],seed[374],seed[767],seed[2180],seed[3302],seed[2154],seed[3383],seed[2492],seed[1956],seed[3765],seed[2350],seed[1636],seed[1120],seed[2569],seed[1158],seed[3023],seed[2191],seed[3283],seed[1804],seed[428],seed[2201],seed[99],seed[2357],seed[2160],seed[334],seed[595],seed[2220],seed[744],seed[1619],seed[1564],seed[1812],seed[3452],seed[1630],seed[2915],seed[3946],seed[673],seed[1385],seed[34],seed[3798],seed[3263],seed[1575],seed[1710],seed[3645],seed[276],seed[1621],seed[1586],seed[1346],seed[3197],seed[2612],seed[1498],seed[2441],seed[3555],seed[3221],seed[3997],seed[477],seed[4023],seed[541],seed[3323],seed[2375],seed[2639],seed[139],seed[494],seed[2885],seed[293],seed[289],seed[15],seed[308],seed[1416],seed[3080],seed[1430],seed[3615],seed[3518],seed[1040],seed[4016],seed[774],seed[1946],seed[2358],seed[1577],seed[3472],seed[436],seed[3698],seed[2836],seed[2165],seed[706],seed[3753],seed[1965],seed[2410],seed[3243],seed[1055],seed[198],seed[913],seed[1478],seed[2643],seed[2944],seed[419],seed[1411],seed[300],seed[1261],seed[1283],seed[3443],seed[3462],seed[3202],seed[2851],seed[347],seed[345],seed[349],seed[97],seed[3205],seed[938],seed[565],seed[917],seed[3773],seed[3007],seed[3703],seed[439],seed[961],seed[825],seed[2509],seed[634],seed[1211],seed[3870],seed[1641],seed[1399],seed[3661],seed[2284],seed[1179],seed[1650],seed[1700],seed[3078],seed[3193],seed[112],seed[1573],seed[286],seed[1721],seed[3606],seed[3421],seed[2234],seed[546],seed[3460],seed[987],seed[3260],seed[1018],seed[2032],seed[2435],seed[170],seed[986],seed[2235],seed[2552],seed[29],seed[2545],seed[960],seed[3459],seed[755],seed[3087],seed[1495],seed[2222],seed[2605],seed[2421],seed[1594],seed[2468],seed[2080],seed[3716],seed[1872],seed[2186],seed[1557],seed[2788],seed[2933],seed[1068],seed[4035],seed[3312],seed[3086],seed[1724],seed[1599],seed[2306],seed[2214],seed[2777],seed[3228],seed[4038],seed[3458],seed[1123],seed[1095],seed[1596],seed[3795],seed[1364],seed[2487],seed[187],seed[1972],seed[2558],seed[711],seed[1470],seed[3829],seed[3764],seed[2957],seed[1080],seed[1923],seed[1589],seed[3804],seed[324],seed[3185],seed[3718],seed[95],seed[1868],seed[2107],seed[1419],seed[1674],seed[1300],seed[1004],seed[1581],seed[3101],seed[839],seed[2990],seed[653],seed[645],seed[3182],seed[3761],seed[2572],seed[3585],seed[3229],seed[3042],seed[3527],seed[1108],seed[1983],seed[3904],seed[823],seed[2582],seed[1013],seed[3238],seed[137],seed[1065],seed[2919],seed[2900],seed[1037],seed[2613],seed[1370],seed[2283],seed[3885],seed[1447],seed[3399],seed[39],seed[1864],seed[2678],seed[3146],seed[1522],seed[2017],seed[3406],seed[415],seed[1808],seed[2633],seed[3583],seed[967],seed[2984],seed[643],seed[3183],seed[480],seed[1827],seed[184],seed[2322],seed[521],seed[786],seed[166],seed[2698],seed[1171],seed[1047],seed[140],seed[806],seed[3571],seed[3580],seed[3563],seed[867],seed[822],seed[805],seed[3621],seed[445],seed[94],seed[3247],seed[1814],seed[4048],seed[2511],seed[553],seed[1747],seed[1566],seed[2708],seed[604],seed[719],seed[281],seed[2039],seed[3649],seed[743],seed[3608],seed[96],seed[1006],seed[3382],seed[955],seed[2942],seed[1221],seed[3572],seed[3329],seed[664],seed[1228],seed[2452],seed[3846],seed[979],seed[3179],seed[3364],seed[3573],seed[2716],seed[637],seed[3415],seed[3110],seed[3426],seed[1350],seed[2528],seed[2127],seed[1775],seed[513],seed[2955],seed[1295],seed[2315],seed[1136],seed[3651],seed[599],seed[333],seed[2460],seed[3512],seed[3944],seed[266],seed[2062],seed[1785],seed[3551],seed[3136],seed[3547],seed[739],seed[1154],seed[1819],seed[3858],seed[1395],seed[2249],seed[3430],seed[2018],seed[3498],seed[537],seed[343],seed[2455],seed[110],seed[3257],seed[1507],seed[752],seed[1223],seed[283],seed[3386],seed[570],seed[3046],seed[1094],seed[113],seed[2610],seed[48],seed[3036],seed[1097],seed[4081],seed[1779],seed[219],seed[159],seed[709],seed[614],seed[197],seed[3950],seed[459],seed[2513],seed[1436],seed[1125],seed[2399],seed[3447],seed[3843],seed[782],seed[4093],seed[3519],seed[3490],seed[688],seed[925],seed[2820],seed[296],seed[3564],seed[3734],seed[3126],seed[1656],seed[1818],seed[731],seed[1948],seed[2373],seed[215],seed[3745],seed[1473],seed[1101],seed[1562],seed[2109],seed[282],seed[393],seed[540],seed[127],seed[2446],seed[695],seed[305],seed[179],seed[3513],seed[4094],seed[2614],seed[956],seed[770],seed[707],seed[2868],seed[3032],seed[71],seed[227],seed[3670],seed[4039],seed[3987],seed[1458],seed[1384],seed[2638],seed[1335],seed[1375],seed[1086],seed[922],seed[2083],seed[980],seed[4014],seed[847],seed[1130],seed[727],seed[2518],seed[1160],seed[560],seed[682],seed[2324],seed[2641],seed[2674],seed[3043],seed[202],seed[3190],seed[3867],seed[3181],seed[2161],seed[3546],seed[3710],seed[524],seed[2556],seed[57],seed[322],seed[621],seed[687],seed[152],seed[2454],seed[532],seed[2884],seed[405],seed[3967],seed[2524],seed[3216],seed[2116],seed[2726],seed[2824],seed[3511],seed[3799],seed[2337],seed[1438],seed[697],seed[2298],seed[3626],seed[3166],seed[1993],seed[2893],seed[1944],seed[1746],seed[88],seed[3326],seed[3533],seed[3791],seed[203],seed[1639],seed[3403],seed[3771],seed[2078],seed[2385],seed[907],seed[3741],seed[1634],seed[603],seed[1561],seed[3892],seed[3909],seed[2684],seed[2765],seed[2309],seed[3900],seed[3966],seed[3969],seed[904],seed[2445],seed[3516],seed[2095],seed[2855],seed[370],seed[273],seed[69],seed[3008],seed[627],seed[1678],seed[58],seed[3424],seed[3816],seed[1272],seed[3053],seed[3196],seed[3448],seed[1609],seed[800],seed[4075],seed[37],seed[2546],seed[2147],seed[2611],seed[2169],seed[2669],seed[3011],seed[3542],seed[2826],seed[2226],seed[3337],seed[1181],seed[2579],seed[2246],seed[1958],seed[3108],seed[3535],seed[1604],seed[3148],seed[1802],seed[587],seed[3747],seed[406],seed[2029],seed[396],seed[3917],seed[1359],seed[1140],seed[1772],seed[2327],seed[2002],seed[2898],seed[932],seed[4092],seed[2805],seed[1099],seed[3543],seed[3310],seed[3971],seed[1041],seed[1007],seed[1688],seed[2263],seed[788],seed[2216],seed[1654],seed[1050],seed[1754],seed[1813],seed[3926],seed[757],seed[16],seed[3015],seed[1889],seed[4070],seed[2535],seed[3418],seed[2767],seed[2368],seed[720],seed[3481],seed[2461],seed[2624],seed[644],seed[3951],seed[353],seed[3276],seed[3203],seed[1111],seed[954],seed[1588],seed[2750],seed[849],seed[155],seed[1787],seed[3290],seed[3920],seed[773],seed[886],seed[2408],seed[4000],seed[2000],seed[1544],seed[1720],seed[1782],seed[394],seed[3125],seed[3135],seed[2929],seed[1028],seed[2849],seed[3150],seed[2432],seed[680],seed[1803],seed[3812],seed[646],seed[3133],seed[465],seed[3206],seed[3976],seed[3392],seed[3685],seed[1658],seed[3152],seed[316],seed[117],seed[765],seed[3120],seed[1301],seed[2051],seed[2390],seed[1343],seed[3865],seed[725],seed[635],seed[3746],seed[3781],seed[1360],seed[2632],seed[2317],seed[2954],seed[3541],seed[591],seed[3888],seed[1026],seed[2903],seed[3278],seed[3737],seed[1199],seed[3497],seed[1468],seed[1693],seed[2046],seed[2227],seed[2706],seed[1250],seed[175],seed[4005],seed[2334],seed[3834],seed[136],seed[3841],seed[3666],seed[3161],seed[4024],seed[45],seed[3173],seed[2371],seed[1928],seed[947],seed[2574],seed[2052],seed[1711],seed[2065],seed[1462],seed[25],seed[1809],seed[3908],seed[2694],seed[3001],seed[3154],seed[2187],seed[1886],seed[368],seed[70],seed[2037],seed[2869],seed[659],seed[1059],seed[1955],seed[2772],seed[1729],seed[1922],seed[462],seed[180],seed[3013],seed[79],seed[3688],seed[2619],seed[3923],seed[1962],seed[3127],seed[2449],seed[2300],seed[3464],seed[2829],seed[3995],seed[3998],seed[1546],seed[3251],seed[331],seed[2500],seed[1051],seed[3780],seed[2850],seed[2508],seed[2704],seed[1119],seed[3832],seed[3111],seed[3823],seed[1551],seed[261],seed[86],seed[2402],seed[3249],seed[2600],seed[2031],seed[3599],seed[1163],seed[995],seed[1264],seed[506],seed[1309],seed[3171],seed[1472],seed[1776],seed[2104],seed[2753],seed[2437],seed[2666],seed[2296],seed[130],seed[2774],seed[2809],seed[1622],seed[3316],seed[1502],seed[1057],seed[1857],seed[172],seed[2677],seed[3974],seed[835],seed[3186],seed[1690],seed[3931],seed[789],seed[1159],seed[12],seed[2681],seed[2909],seed[2662],seed[2622],seed[1837],seed[2172],seed[2895],seed[1252],seed[2737],seed[3943],seed[1714],seed[2961],seed[3544],seed[3863],seed[3393],seed[3217],seed[1241],seed[1815],seed[3062],seed[2013],seed[654],seed[2691],seed[3066],seed[3455],seed[1701],seed[1345],seed[31],seed[3930],seed[2325],seed[89],seed[1835],seed[2872],seed[3553],seed[488],seed[1517],seed[3461],seed[2444],seed[3239],seed[2649],seed[509],seed[2336],seed[2310],seed[373],seed[2431],seed[1696],seed[2739],seed[3751],seed[2418],seed[3277],seed[461],seed[3906],seed[2276],seed[3866],seed[3451],seed[1293],seed[2070],seed[3242],seed[173],seed[1512],seed[1249],seed[1524],seed[3794],seed[3099],seed[683],seed[2858],seed[733],seed[1227],seed[3646],seed[417],seed[1011],seed[3857],seed[3524],seed[670],seed[103],seed[2028],seed[4030],seed[407],seed[574],seed[46],seed[2190],seed[2979],seed[819],seed[290],seed[2997],seed[4032],seed[1190],seed[1832],seed[3595],seed[195],seed[3935],seed[821],seed[978],seed[83],seed[2166],seed[1195],seed[3956],seed[2185],seed[2079],seed[3522],seed[704],seed[142],seed[615],seed[1187],seed[1892],seed[2286],seed[2288],seed[3140],seed[1009],seed[1734],seed[3289],seed[47],seed[816],seed[1319],seed[3293],seed[3348],seed[366],seed[400],seed[2364],seed[3709],seed[1117],seed[1774],seed[210],seed[1821],seed[2950],seed[1424],seed[2804],seed[2091],seed[185],seed[44],seed[342],seed[129],seed[1316],seed[3003],seed[3782],seed[1628],seed[2761],seed[3830],seed[3049],seed[3371],seed[3984],seed[1387],seed[2617],seed[539],seed[1705],seed[49],seed[3788],seed[2010],seed[2040],seed[1204],seed[3355],seed[2429],seed[794],seed[3752],seed[3407],seed[1302],seed[1471],seed[2277],seed[199],seed[171],seed[1292],seed[1651],seed[1558],seed[1475],seed[2030],seed[3662],seed[3338],seed[916],seed[3778],seed[1398],seed[2114],seed[935],seed[3730],seed[1185],seed[675],seed[2099],seed[397],seed[272],seed[1552],seed[2542],seed[2779],seed[3985],seed[582],seed[2891],seed[2635],seed[2519],seed[3031],seed[2274],seed[440],seed[581],seed[2285],seed[3558],seed[703],seed[1924],seed[1153],seed[2626],seed[921],seed[1968],seed[2121],seed[2789],seed[2174],seed[3419],seed[1875],seed[327],seed[317],seed[3391],seed[2601],seed[3978],seed[802],seed[1365],seed[912],seed[2887],seed[4037],seed[3330],seed[2964],seed[1450],seed[377],seed[220],seed[1021],seed[1511],seed[3105],seed[3992],seed[3219],seed[2486],seed[1602],seed[1353],seed[128],seed[4006],seed[1349],seed[2178],seed[325],seed[642],seed[678],seed[690],seed[3332],seed[11],seed[454],seed[1740],seed[3076],seed[716],seed[629],seed[2205],seed[3561],seed[3294],seed[1382],seed[161],seed[3559],seed[1180],seed[153],seed[1769],seed[1344],seed[367],seed[1743],seed[3972],seed[2770],seed[43],seed[1598],seed[339],seed[571],seed[2864],seed[1554],seed[557],seed[1597],seed[1129],seed[1445],seed[1407],seed[3845],seed[2948],seed[1662],seed[1453],seed[3162],seed[3093],seed[1166],seed[2311],seed[2250],seed[1242],seed[93],seed[475],seed[2261],seed[292],seed[803],seed[255],seed[4002],seed[2875],seed[2660],seed[1107],seed[1217],seed[2575],seed[2935],seed[3040],seed[2025],seed[3854],seed[1735],seed[2360],seed[829],seed[229],seed[1781],seed[3844],seed[1854],seed[2963],seed[7],seed[1031],seed[699],seed[1491],seed[993],seed[846],seed[211],seed[87],seed[1352],seed[1777],seed[3299],seed[205],seed[2329],seed[2515],seed[734],seed[1679],seed[2491],seed[3137],seed[2221],seed[3648],seed[3569],seed[132],seed[3530],seed[2873],seed[1056],seed[3098],seed[2842],seed[3097],seed[3570],seed[768],seed[1192],seed[742],seed[2370],seed[1974],seed[3204],seed[2966],seed[158],seed[1971],seed[1333],seed[1061],seed[647],seed[2897],seed[3625],seed[2458],seed[297],seed[3665],seed[1992],seed[2346],seed[3942],seed[738],seed[3489],seed[2987],seed[2347],seed[1276],seed[3441],seed[1778],seed[3676],seed[495],seed[545],seed[3083],seed[1046],seed[2917],seed[254],seed[2457],seed[968],seed[1500],seed[889],seed[997],seed[556],seed[1053],seed[2507],seed[606],seed[2553],seed[2450],seed[3390],seed[3818],seed[785],seed[2688],seed[3057],seed[3212],seed[1712],seed[1885],seed[962],seed[4034],seed[2326],seed[3777],seed[3039],seed[975],seed[2938],seed[2240],seed[3770],seed[2237],seed[2985],seed[2430],seed[3678],seed[3096],seed[2003],seed[2170],seed[357],seed[3054],seed[2644],seed[1840],seed[2453],seed[3723],seed[3952],seed[3576],seed[2481],seed[4063],seed[1446],seed[1532],seed[1210],seed[2314],seed[3139],seed[303],seed[2269],seed[1984],seed[1168],seed[62],seed[403],seed[1506],seed[3839],seed[2202],seed[717],seed[3144],seed[4065],seed[1685],seed[1320],seed[1670],seed[2392],seed[3958],seed[3158],seed[1811],seed[860],seed[3957],seed[2268],seed[13],seed[133],seed[3104],seed[686],seed[3915],seed[222],seed[3597],seed[2778],seed[2094],seed[853],seed[213],seed[977],seed[3091],seed[708],seed[3496],seed[1245],seed[3528],seed[758],seed[3617],seed[2252],seed[1726],seed[1518],seed[3640],seed[2760],seed[4079],seed[3581],seed[3815],seed[3450],seed[8],seed[1172],seed[468],seed[976],seed[1988],seed[1298],seed[1994],seed[498],seed[332],seed[3408],seed[1866],seed[879],seed[90],seed[3288],seed[2506],seed[1452],seed[1404],seed[1257],seed[3514],seed[2442],seed[2970],seed[861],seed[2182],seed[1202],seed[2379],seed[64],seed[1605],seed[2892],seed[596],seed[840],seed[592],seed[520],seed[1969],seed[651],seed[3949],seed[3187],seed[3255],seed[899],seed[399],seed[2673],seed[1282],seed[1541],seed[1147],seed[630],seed[1176],seed[2102],seed[115],seed[1089],seed[1493],seed[1680],seed[3766],seed[1805],seed[2798],seed[1441],seed[2802],seed[3331],seed[2562],seed[256],seed[1016],seed[3993],seed[3306],seed[942],seed[3921],seed[2797],seed[3339],seed[931],seed[2874],seed[100],seed[3044],seed[684],seed[2862],seed[1036],seed[2854],seed[1616],seed[2571],seed[2297],seed[3653],seed[929],seed[3848],seed[3954],seed[302],seed[2597],seed[1917],seed[2537],seed[1728],seed[275],seed[249],seed[2264],seed[575],seed[723],seed[463],seed[1014],seed[1613],seed[844],seed[1290],seed[1278],seed[756],seed[2847],seed[1698],seed[2819],seed[3484],seed[188],seed[59],seed[623],seed[3079],seed[3862],seed[2936],seed[1480],seed[2301],seed[3285],seed[2072],seed[244],seed[3690],seed[984],seed[3010],seed[2616],seed[1066],seed[722],seed[3357],seed[1836],seed[453],seed[3824],seed[1337],seed[2257],seed[928],seed[3894],seed[3775],seed[1164],seed[2006],seed[1281],seed[1768],seed[3412],seed[3929],seed[3801],seed[2714],seed[1306],seed[2700],seed[3864],seed[1487],seed[2563],seed[3258],seed[1391],seed[2870],seed[3902],seed[1076],seed[779],seed[125],seed[554],seed[2960],seed[1881],seed[666],seed[1989],seed[2830],seed[945],seed[455],seed[2490],seed[988],seed[2480],seed[2712],seed[2766],seed[1888],seed[1448],seed[3790],seed[2554],seed[1862],seed[2464],seed[437],seed[609],seed[1128],seed[2776],seed[1861],seed[3072],seed[941],seed[2530],seed[2534],seed[837],seed[1741],seed[910],seed[1527],seed[648],seed[3377],seed[299],seed[1386],seed[663],seed[395],seed[2682],seed[3711],seed[2426],seed[1331],seed[4010],seed[108],seed[3808],seed[2692],seed[3232],seed[3634],seed[625],seed[1167],seed[1607],seed[3849],seed[3601],seed[2241],seed[1173],seed[3609],seed[1786],seed[3164],seed[2145],seed[3627],seed[398],seed[3655],seed[3600],seed[2231],seed[3423],seed[2332],seed[3246],seed[969],seed[1833],seed[1788],seed[1012],seed[239],seed[401],seed[3567],seed[1113],seed[843],seed[583],seed[926],seed[1576],seed[3463],seed[1025],seed[1987],seed[3414],seed[3629],seed[2670],seed[875],seed[3814],seed[4090],seed[2756],seed[1],seed[2585],seed[3717],seed[2427],seed[3523],seed[2389],seed[572],seed[2646],seed[2292],seed[2338],seed[238],seed[217],seed[2578],seed[4019],seed[877],seed[512],seed[1841],seed[1846],seed[2588],seed[1933],seed[965],seed[2401],seed[1790],seed[156],seed[1085],seed[3132],seed[2016],seed[486],seed[2484],seed[1816],seed[2713],seed[510],seed[427],seed[3284],seed[2980],seed[2496],seed[3568],seed[3029],seed[1896],seed[1996],seed[2541],seed[972],seed[2438],seed[1400],seed[3560],seed[1356],seed[1759],seed[801],seed[2520],seed[3591],seed[3647],seed[3473],seed[2952],seed[679],seed[2566],seed[1481],seed[3400],seed[892],seed[2881],seed[2020],seed[3874],seed[1555],seed[1727],seed[77],seed[1401],seed[193],seed[3347],seed[3669],seed[4020],seed[201],seed[1488],seed[2672],seed[1460],seed[668],seed[3619],seed[534],seed[598],seed[3177],seed[602],seed[1751],seed[1839],seed[718],seed[3273],seed[2699],seed[1758],seed[2655],seed[1437],seed[2642],seed[2258],seed[2118],seed[2412],seed[288],seed[4036],seed[890],seed[3611],seed[1288],seed[4047],seed[1838],seed[3840],seed[3499],seed[2941],seed[1547],seed[1947],seed[1482],seed[597],seed[147],seed[2501],seed[2063],seed[3075],seed[3719],seed[3507],seed[2799],seed[1048],seed[154],seed[842],seed[2290],seed[3733],seed[754],seed[3534],seed[2203],seed[970],seed[3953],seed[364],seed[307],seed[501],seed[3859],seed[2248],seed[4057],seed[3725],seed[2398],seed[1467],seed[269],seed[3081],seed[1403],seed[186],seed[2448],seed[176],seed[432],seed[2047],seed[3936],seed[2793],seed[836],seed[1767],seed[824],seed[2573],seed[1697],seed[1870],seed[966],seed[233],seed[375],seed[423],seed[2735],seed[1528],seed[2215],seed[2911],seed[2092],seed[661],seed[1358],seed[1138],seed[3379],seed[2343],seed[150],seed[2108],seed[429],seed[386],seed[2469],seed[2806],seed[3736],seed[671],seed[1069],seed[3650],seed[1000],seed[1501],seed[3783],seed[2024],seed[3509],seed[1311],seed[2112],seed[1671],seed[433],seed[123],seed[2305],seed[1504],seed[3385],seed[3396],seed[710],seed[2920],seed[2992],seed[3397],seed[3721],seed[2238],seed[1663],seed[891],seed[2514],seed[3982],seed[2397],seed[2974],seed[335],seed[1752],seed[3027],seed[3707],seed[2512],seed[2244],seed[2321],seed[2245],seed[2640],seed[628],seed[2932],seed[2333],seed[4033],seed[1629],seed[3266],seed[881],seed[497],seed[3769],seed[2113],seed[4058],seed[730],seed[2105],seed[1521],seed[3973],seed[3114],seed[3940],seed[1499],seed[3644],seed[3267],seed[3109],seed[1939],seed[3292],seed[387],seed[51],seed[2539],seed[3056],seed[3979],seed[612],seed[2228],seed[746],seed[3103],seed[3545],seed[3313],seed[2757],seed[3262],seed[75],seed[2822],seed[3005],seed[4066],seed[221],seed[721],seed[1112],seed[385],seed[769],seed[1357],seed[530],seed[493],seed[1640],seed[3123],seed[3510],seed[2097],seed[2982],seed[3404],seed[2607],seed[2383],seed[3026],seed[3557],seed[1736],seed[3726],seed[2377],seed[992],seed[735],seed[1748],seed[3880],seed[1925],seed[2156],seed[3456],seed[3089],seed[2594],seed[652],seed[2721],seed[1953],seed[1514],seed[2695],seed[2719],seed[2593],seed[3082],seed[1667],seed[2417],seed[3287],seed[3875],seed[1332],seed[2843],seed[1289],seed[1990],seed[1973],seed[1920],seed[845],seed[1657],seed[2910],seed[1945],seed[2618],seed[2403],seed[435],seed[3700],seed[566],seed[1677],seed[1709],seed[1392],seed[792],seed[2595],seed[2631],seed[204],seed[1592],seed[3130],seed[1201],seed[2926],seed[3160],seed[182],seed[4025],seed[1121],seed[2061],seed[3789],seed[3004],seed[1686],seed[450],seed[1200],seed[3637],seed[2785],seed[340],seed[3025],seed[1676],seed[1247],seed[1959],seed[3827],seed[3884],seed[2548],seed[2106],seed[1265],seed[1443],seed[2451],seed[228],seed[42],seed[2705],seed[3058],seed[3668],seed[3856],seed[3501],seed[1203],seed[2840],seed[27],seed[2271],seed[827],seed[1545],seed[525],seed[2598],seed[2922],seed[1660],seed[1023],seed[865],seed[3134],seed[209],seed[2560],seed[3014],seed[346],seed[3633],seed[3587],seed[1921],seed[1764],seed[641],seed[3879],seed[2683],seed[1409],seed[3131],seed[3409],seed[2082],seed[3349],seed[1673],seed[1887],seed[2318],seed[2175],seed[251],seed[3860],seed[1543],seed[379],seed[1444],seed[3195],seed[1580],seed[2775],seed[2055],seed[3842],seed[1624],seed[2151],seed[2242],seed[313],seed[1600],seed[936],seed[894],seed[3642],seed[250],seed[852],seed[200],seed[3318],seed[2734],seed[2144],seed[3437],seed[1474],seed[2320],seed[2953],seed[833],seed[2436],seed[2801],seed[1137],seed[818],seed[905],seed[56],seed[2902],seed[1383],seed[443],seed[3889],seed[3887],seed[2413],seed[2504],seed[1716],seed[1362],seed[2090],seed[1131],seed[3566],seed[1496],seed[1903],seed[2213],seed[2117],seed[280],seed[952],seed[1873],seed[3315],seed[3614],seed[2341],seed[3333],seed[323],seed[1824],seed[3107],seed[2879],seed[2362],seed[2581],seed[2732],seed[3831],seed[2189],seed[2880],seed[1145],seed[1858],seed[2064],seed[2833],seed[2736],seed[1961],seed[4071],seed[1406],seed[2702],seed[298],seed[2584],seed[2393],seed[491],seed[1603],seed[2939],seed[1916],seed[3910],seed[1104],seed[2807],seed[3999],seed[3055],seed[624],seed[543],seed[750],seed[1906],seed[1189],seed[2993],seed[2084],seed[1237],seed[2351],seed[3632],seed[2967],seed[1898],seed[2372],seed[264],seed[2304],seed[3446],seed[2168],seed[1428],seed[2628],seed[2056],seed[3395],seed[3192],seed[964],seed[1516],seed[2589],seed[3549],seed[1717],seed[3256],seed[3712],seed[1479],seed[866],seed[3298],seed[356],seed[1523],seed[2008],seed[360],seed[1584],seed[862],seed[1230],seed[2229],seed[235],seed[206],seed[2853],seed[2353],seed[3453],seed[4054],seed[3465],seed[2591],seed[1188],seed[3853],seed[3502],seed[3590],seed[1170],seed[1234],seed[1952],seed[1538],seed[527],seed[478],seed[2243],seed[3122],seed[729],seed[1649],seed[3835],seed[4089],seed[3362],seed[2791],seed[1723],seed[354],seed[640],seed[3699],seed[2889],seed[3328],seed[194],seed[3714],seed[1027],seed[2289],seed[590],seed[3454],seed[30],seed[1978],seed[1559],seed[3270],seed[21],seed[2081],seed[1116],seed[3153],seed[656],seed[605],seed[1141],seed[1148],seed[1127],seed[177],seed[2821],seed[728],seed[2841],seed[2894],seed[2969],seed[4045],seed[3064],seed[3170],seed[1851],seed[1975],seed[622],seed[3468],seed[3988],seed[2485],seed[212],seed[2192],seed[4056],seed[3245],seed[2044],seed[3100],seed[2679],seed[3281],seed[1035],seed[2054],seed[2568],seed[1156],seed[4004],seed[3225],seed[1100],seed[3540],seed[1606],seed[1142],seed[1757],seed[3358],seed[1212],seed[1761],seed[2312],seed[330],seed[3941],seed[3359],seed[4060],seed[3033],seed[751],seed[473],seed[3602],seed[111],seed[1612],seed[943],seed[1033],seed[3405],seed[3945],seed[3340],seed[2857],seed[883],seed[1280],seed[3613],seed[3525],seed[474],seed[639],seed[780],seed[2022],seed[691],seed[713],seed[3607],seed[3592],seed[1849],seed[2718],seed[1461],seed[2690],seed[1668],seed[511],seed[3469],seed[178],seed[3715],seed[1231],seed[1347],seed[1291],seed[813],seed[3792],seed[311],seed[2752],seed[3002],seed[793],seed[3720],seed[3521],seed[3492],seed[3822],seed[3065],seed[1661],seed[1810],seed[3833],seed[3873],seed[2972],seed[3275],seed[3656],seed[901],seed[2828],seed[3020],seed[2302],seed[3048],seed[3435],seed[4027],seed[3483],seed[138],seed[608],seed[617],seed[2965],seed[3209],seed[2380],seed[1177],seed[1807],seed[4091],seed[2918],seed[2466],seed[3494],seed[884],seed[1198],seed[1937],seed[14],seed[3411],seed[3691],seed[3526],seed[4087],seed[1312],seed[109],seed[1115],seed[1422],seed[1328],seed[1733],seed[421],seed[2609],seed[1852],seed[3006],seed[2462],seed[1763],seed[216],seed[61],seed[2021],seed[1542],seed[82],seed[2923],seed[2253],seed[1477],seed[337],seed[3102],seed[858],seed[2382],seed[1476],seed[1863],seed[1665],seed[576],seed[2291],seed[3342],seed[2313],seed[1871],seed[3045],seed[855],seed[1550],seed[2818],seed[3157],seed[267],seed[3628],seed[3838],seed[1715],seed[3180],seed[508],seed[2255],seed[3308]}),
        .cross_prob(cross_prob),
        .codeword(codeword9),
        .received(received9)
        );
    
    bsc bsc10(
        .clk(clk),
        .reset(reset),
        .seed({seed[3624],seed[2102],seed[1027],seed[2471],seed[3952],seed[3977],seed[2390],seed[521],seed[611],seed[1731],seed[624],seed[2913],seed[990],seed[1577],seed[3172],seed[80],seed[3010],seed[2263],seed[793],seed[582],seed[2671],seed[3186],seed[1654],seed[2864],seed[199],seed[3321],seed[1964],seed[3311],seed[1230],seed[4060],seed[1850],seed[3641],seed[2979],seed[2823],seed[1375],seed[4041],seed[699],seed[3877],seed[1942],seed[2009],seed[3599],seed[457],seed[1921],seed[3659],seed[2425],seed[3963],seed[2162],seed[861],seed[2616],seed[2987],seed[3047],seed[2444],seed[3861],seed[325],seed[2833],seed[3203],seed[2954],seed[671],seed[1005],seed[2686],seed[112],seed[2034],seed[1420],seed[753],seed[3388],seed[1327],seed[89],seed[202],seed[777],seed[1208],seed[2882],seed[4065],seed[353],seed[2972],seed[1885],seed[190],seed[3],seed[3727],seed[1744],seed[1745],seed[885],seed[77],seed[1185],seed[1038],seed[2600],seed[887],seed[2801],seed[3718],seed[3444],seed[2218],seed[529],seed[680],seed[1879],seed[4066],seed[967],seed[3291],seed[40],seed[3192],seed[3643],seed[238],seed[2769],seed[2052],seed[2473],seed[1514],seed[1310],seed[2347],seed[3269],seed[1968],seed[2876],seed[2412],seed[1549],seed[2664],seed[1379],seed[3839],seed[808],seed[2803],seed[2003],seed[2295],seed[1993],seed[1155],seed[550],seed[700],seed[1334],seed[3306],seed[3316],seed[1153],seed[1837],seed[2525],seed[713],seed[2441],seed[1352],seed[729],seed[64],seed[348],seed[1887],seed[2970],seed[595],seed[3805],seed[1688],seed[870],seed[1233],seed[1878],seed[368],seed[3993],seed[419],seed[4074],seed[274],seed[2279],seed[1930],seed[3268],seed[203],seed[2842],seed[3240],seed[1010],seed[1068],seed[2812],seed[2495],seed[1637],seed[2649],seed[1796],seed[3767],seed[2507],seed[1540],seed[3348],seed[590],seed[2024],seed[3602],seed[50],seed[3353],seed[1762],seed[1965],seed[2221],seed[2054],seed[342],seed[3800],seed[207],seed[2593],seed[1316],seed[3809],seed[1623],seed[6],seed[286],seed[344],seed[2381],seed[3079],seed[1210],seed[2017],seed[1291],seed[302],seed[1363],seed[946],seed[1950],seed[3214],seed[2504],seed[4087],seed[1618],seed[2108],seed[3420],seed[997],seed[371],seed[1365],seed[2258],seed[2070],seed[2701],seed[952],seed[129],seed[2008],seed[3006],seed[16],seed[244],seed[1324],seed[553],seed[3096],seed[367],seed[2318],seed[2532],seed[1227],seed[3329],seed[2627],seed[1404],seed[3971],seed[1614],seed[4059],seed[1458],seed[685],seed[375],seed[3464],seed[1919],seed[2125],seed[2084],seed[773],seed[3666],seed[3127],seed[597],seed[2016],seed[575],seed[1653],seed[1364],seed[1643],seed[489],seed[3499],seed[1106],seed[642],seed[1561],seed[1438],seed[470],seed[18],seed[1289],seed[733],seed[1518],seed[2528],seed[97],seed[544],seed[663],seed[3537],seed[4075],seed[669],seed[1882],seed[3675],seed[3867],seed[888],seed[3872],seed[1550],seed[2937],seed[2784],seed[2486],seed[219],seed[2524],seed[641],seed[31],seed[113],seed[3454],seed[2587],seed[1719],seed[1773],seed[2406],seed[3121],seed[963],seed[1441],seed[973],seed[2091],seed[3290],seed[3275],seed[235],seed[2929],seed[3583],seed[3597],seed[100],seed[2834],seed[3563],seed[2130],seed[2362],seed[2297],seed[2619],seed[1860],seed[3983],seed[2517],seed[3086],seed[467],seed[288],seed[1865],seed[4002],seed[3802],seed[2632],seed[2777],seed[155],seed[3526],seed[3038],seed[622],seed[2299],seed[762],seed[2974],seed[532],seed[1689],seed[1813],seed[410],seed[2774],seed[2867],seed[2621],seed[159],seed[3202],seed[1279],seed[2339],seed[3961],seed[1533],seed[3535],seed[1362],seed[229],seed[1013],seed[4022],seed[554],seed[2180],seed[1666],seed[1682],seed[95],seed[2199],seed[991],seed[123],seed[989],seed[1201],seed[676],seed[471],seed[56],seed[662],seed[3950],seed[1408],seed[1048],seed[1202],seed[29],seed[2531],seed[3881],seed[2661],seed[1353],seed[2436],seed[1923],seed[3387],seed[2958],seed[3527],seed[2626],seed[1121],seed[3441],seed[3572],seed[1248],seed[2107],seed[2004],seed[1803],seed[3377],seed[795],seed[2453],seed[4037],seed[2167],seed[2551],seed[605],seed[694],seed[1394],seed[3492],seed[2676],seed[2918],seed[1284],seed[1736],seed[2432],seed[3631],seed[1576],seed[1782],seed[679],seed[1189],seed[2113],seed[2442],seed[42],seed[486],seed[3895],seed[668],seed[2350],seed[3391],seed[376],seed[2560],seed[1077],seed[2602],seed[1494],seed[3813],seed[1465],seed[426],seed[3147],seed[2206],seed[4025],seed[3264],seed[2492],seed[3518],seed[717],seed[591],seed[2811],seed[160],seed[3515],seed[3789],seed[3978],seed[2591],seed[3610],seed[2831],seed[3236],seed[53],seed[407],seed[381],seed[339],seed[301],seed[3178],seed[953],seed[839],seed[90],seed[1396],seed[3762],seed[3663],seed[2853],seed[581],seed[1370],seed[552],seed[1390],seed[1181],seed[3614],seed[4033],seed[1239],seed[2150],seed[2076],seed[1672],seed[1466],seed[3893],seed[828],seed[2756],seed[2706],seed[652],seed[646],seed[2251],seed[1815],seed[1109],seed[3764],seed[2051],seed[2730],seed[3029],seed[3892],seed[1099],seed[1145],seed[38],seed[2977],seed[718],seed[2982],seed[3953],seed[1501],seed[1816],seed[1806],seed[4034],seed[2061],seed[3104],seed[7],seed[386],seed[2173],seed[8],seed[945],seed[3401],seed[2553],seed[3714],seed[1909],seed[838],seed[1776],seed[3976],seed[3871],seed[2338],seed[3836],seed[1510],seed[1044],seed[2767],seed[1366],seed[3386],seed[380],seed[1030],seed[1384],seed[720],seed[3513],seed[485],seed[3141],seed[3865],seed[3123],seed[2343],seed[3365],seed[2422],seed[2168],seed[2097],seed[2681],seed[2566],seed[3347],seed[3342],seed[304],seed[2576],seed[3571],seed[922],seed[1599],seed[3003],seed[2790],seed[3285],seed[3379],seed[1344],seed[3848],seed[2736],seed[2185],seed[1624],seed[2021],seed[2922],seed[3191],seed[834],seed[1183],seed[3668],seed[2376],seed[2465],seed[1073],seed[3734],seed[3399],seed[1972],seed[3937],seed[975],seed[1276],seed[2253],seed[243],seed[3901],seed[4070],seed[1251],seed[2967],seed[3238],seed[3355],seed[960],seed[4010],seed[142],seed[3906],seed[1931],seed[4067],seed[2928],seed[2691],seed[3065],seed[3448],seed[3325],seed[3590],seed[1246],seed[763],seed[1405],seed[3760],seed[3022],seed[1409],seed[3478],seed[2100],seed[3676],seed[1461],seed[523],seed[463],seed[1709],seed[2605],seed[2244],seed[3480],seed[1794],seed[2692],seed[1301],seed[464],seed[647],seed[545],seed[1308],seed[3930],seed[2386],seed[4021],seed[101],seed[1900],seed[3181],seed[1977],seed[2699],seed[3260],seed[1026],seed[1385],seed[1329],seed[3049],seed[3462],seed[1095],seed[2788],seed[2696],seed[1676],seed[623],seed[1870],seed[2521],seed[3905],seed[854],seed[213],seed[1867],seed[1932],seed[4081],seed[2171],seed[3699],seed[3818],seed[3274],seed[2796],seed[1224],seed[172],seed[1267],seed[2641],seed[3646],seed[1893],seed[2990],seed[1262],seed[2943],seed[109],seed[1785],seed[2237],seed[2188],seed[108],seed[3942],seed[3775],seed[1740],seed[3859],seed[1051],seed[1292],seed[1567],seed[1031],seed[1836],seed[772],seed[3050],seed[1916],seed[2588],seed[2570],seed[1123],seed[3018],seed[1045],seed[287],seed[787],seed[1890],seed[1403],seed[3258],seed[1434],seed[931],seed[3284],seed[2715],seed[2994],seed[200],seed[3541],seed[2538],seed[1430],seed[72],seed[2565],seed[2844],seed[4038],seed[2885],seed[1165],seed[2836],seed[502],seed[59],seed[2154],seed[361],seed[1674],seed[3195],seed[1874],seed[20],seed[2215],seed[1772],seed[744],seed[869],seed[3507],seed[3974],seed[1088],seed[775],seed[3265],seed[1256],seed[2648],seed[1543],seed[188],seed[3918],seed[1767],seed[3402],seed[4077],seed[496],seed[3728],seed[1553],seed[1221],seed[490],seed[1842],seed[3148],seed[3551],seed[3980],seed[3320],seed[192],seed[3736],seed[2326],seed[3570],seed[2233],seed[2888],seed[3432],seed[1895],seed[2625],seed[2035],seed[1187],seed[3054],seed[3281],seed[1573],seed[3725],seed[2332],seed[444],seed[415],seed[688],seed[3594],seed[390],seed[2757],seed[413],seed[3826],seed[1317],seed[3075],seed[3709],seed[2606],seed[2179],seed[425],seed[2980],seed[3481],seed[2157],seed[3294],seed[1941],seed[345],seed[561],seed[1280],seed[892],seed[3058],seed[2117],seed[1053],seed[3987],seed[1186],seed[247],seed[2829],seed[2624],seed[1297],seed[48],seed[166],seed[2282],seed[1075],seed[1512],seed[3163],seed[955],seed[1451],seed[3383],seed[1231],seed[2449],seed[193],seed[312],seed[1036],seed[3595],seed[1961],seed[895],seed[473],seed[3738],seed[2724],seed[3630],seed[1499],seed[3863],seed[2969],seed[248],seed[3740],seed[2945],seed[1278],seed[2557],seed[1046],seed[875],seed[465],seed[2577],seed[1303],seed[249],seed[3791],seed[1617],seed[3864],seed[592],seed[3639],seed[3811],seed[451],seed[3463],seed[3529],seed[3187],seed[3620],seed[1597],seed[2192],seed[827],seed[1305],seed[659],seed[3223],seed[2044],seed[328],seed[3868],seed[3426],seed[3221],seed[958],seed[886],seed[436],seed[2181],seed[3210],seed[3707],seed[804],seed[1949],seed[1454],seed[2055],seed[388],seed[927],seed[252],seed[3785],seed[1701],seed[1537],seed[2516],seed[3549],seed[2629],seed[1655],seed[2095],seed[3522],seed[801],seed[3884],seed[1012],seed[684],seed[537],seed[3622],seed[3917],seed[770],seed[3453],seed[1098],seed[969],seed[3770],seed[3502],seed[3466],seed[2592],seed[2909],seed[3697],seed[693],seed[3504],seed[3889],seed[315],seed[1505],seed[3632],seed[633],seed[2195],seed[2890],seed[3136],seed[3002],seed[1448],seed[515],seed[1875],seed[1360],seed[3082],seed[3514],seed[2445],seed[1866],seed[3810],seed[3312],seed[2018],seed[2333],seed[1832],seed[3609],seed[3354],seed[1605],seed[3640],seed[1631],seed[2825],seed[210],seed[2750],seed[2300],seed[1275],seed[4086],seed[2223],seed[1557],seed[2307],seed[1983],seed[3053],seed[2948],seed[4095],seed[2512],seed[3298],seed[2291],seed[1862],seed[196],seed[1928],seed[867],seed[3324],seed[3220],seed[1716],seed[842],seed[3682],seed[2861],seed[877],seed[133],seed[482],seed[3579],seed[3706],seed[2628],seed[3370],seed[2871],seed[1523],seed[578],seed[3841],seed[2760],seed[3660],seed[1873],seed[769],seed[850],seed[4043],seed[1804],seed[2446],seed[2415],seed[3156],seed[1054],seed[1376],seed[3175],seed[703],seed[802],seed[2371],seed[765],seed[73],seed[3756],seed[69],seed[1489],seed[3858],seed[2367],seed[782],seed[321],seed[3914],seed[3144],seed[2499],seed[385],seed[2615],seed[1180],seed[2776],seed[2995],seed[3479],seed[2418],seed[2510],seed[1864],seed[2865],seed[3201],seed[1955],seed[3211],seed[1049],seed[1651],seed[3512],seed[585],seed[826],seed[1287],seed[2976],seed[640],seed[2848],seed[3543],seed[3036],seed[1978],seed[276],seed[1675],seed[517],seed[2152],seed[593],seed[851],seed[3157],seed[3247],seed[1626],seed[71],seed[2145],seed[768],seed[2459],seed[2014],seed[357],seed[1791],seed[2781],seed[3305],seed[897],seed[3028],seed[2312],seed[3411],seed[796],seed[3188],seed[3866],seed[1001],seed[1673],seed[156],seed[551],seed[3131],seed[3729],seed[2485],seed[1506],seed[2940],seed[3880],seed[2461],seed[300],seed[3951],seed[1632],seed[2753],seed[1940],seed[833],seed[1177],seed[1750],seed[3975],seed[191],seed[3510],seed[1338],seed[1869],seed[1061],seed[1527],seed[2121],seed[2193],seed[1421],seed[2169],seed[3382],seed[2711],seed[2401],seed[3717],seed[2464],seed[2110],seed[686],seed[2610],seed[574],seed[1758],seed[1226],seed[3705],seed[2944],seed[1733],seed[4027],seed[3259],seed[3118],seed[3442],seed[2794],seed[2103],seed[3996],seed[1811],seed[3523],seed[1880],seed[1126],seed[2092],seed[1713],seed[1406],seed[3552],seed[1229],seed[3553],seed[2281],seed[3056],seed[3485],seed[2733],seed[589],seed[2216],seed[3032],seed[2973],seed[3908],seed[813],seed[2346],seed[4045],seed[608],seed[3343],seed[1903],seed[745],seed[1560],seed[2151],seed[2907],seed[1821],seed[3369],seed[3425],seed[2642],seed[3856],seed[2806],seed[1566],seed[3012],seed[3840],seed[131],seed[3278],seed[1070],seed[513],seed[165],seed[1554],seed[1337],seed[1111],seed[268],seed[3698],seed[3431],seed[2132],seed[906],seed[1858],seed[122],seed[752],seed[634],seed[1485],seed[1948],seed[362],seed[476],seed[725],seed[2294],seed[2226],seed[1535],seed[1169],seed[1629],seed[2264],seed[2997],seed[1372],seed[3437],seed[3069],seed[0],seed[1906],seed[3048],seed[1004],seed[130],seed[177],seed[2868],seed[2849],seed[455],seed[1603],seed[577],seed[3174],seed[872],seed[3461],seed[3757],seed[1160],seed[23],seed[3506],seed[3153],seed[1008],seed[222],seed[2562],seed[1288],seed[937],seed[3132],seed[1578],seed[1339],seed[1072],seed[1795],seed[2703],seed[1319],seed[785],seed[1002],seed[3931],seed[3129],seed[1043],seed[1622],seed[3967],seed[2644],seed[4015],seed[4084],seed[125],seed[497],seed[1402],seed[2575],seed[1551],seed[2277],seed[1802],seed[3773],seed[3907],seed[4072],seed[1196],seed[761],seed[2342],seed[63],seed[3860],seed[3081],seed[1151],seed[2447],seed[1516],seed[2093],seed[571],seed[3396],seed[240],seed[259],seed[1924],seed[211],seed[2058],seed[3073],seed[3519],seed[4013],seed[1014],seed[3176],seed[2136],seed[136],seed[1175],seed[1323],seed[3779],seed[127],seed[2454],seed[1315],seed[2534],seed[3687],seed[3517],seed[2859],seed[2306],seed[2941],seed[3703],seed[555],seed[3766],seed[1184],seed[3219],seed[47],seed[2398],seed[1133],seed[3165],seed[2673],seed[3031],seed[184],seed[3629],seed[1140],seed[2419],seed[3286],seed[3711],seed[3801],seed[3429],seed[904],seed[4011],seed[2942],seed[3611],seed[4051],seed[2078],seed[2420],seed[460],seed[2573],seed[331],seed[3684],seed[3405],seed[1558],seed[1055],seed[1582],seed[3322],seed[2259],seed[1393],seed[1742],seed[2334],seed[2988],seed[1741],seed[563],seed[146],seed[212],seed[1593],seed[2275],seed[2187],seed[2545],seed[2252],seed[1640],seed[492],seed[1234],seed[378],seed[1418],seed[1702],seed[54],seed[982],seed[1780],seed[420],seed[1429],seed[3695],seed[3193],seed[560],seed[2402],seed[433],seed[2579],seed[4006],seed[631],seed[1074],seed[458],seed[3566],seed[2348],seed[1225],seed[1926],seed[1824],seed[2175],seed[2205],seed[3057],seed[876],seed[475],seed[2939],seed[3591],seed[1747],seed[1479],seed[1199],seed[1057],seed[3470],seed[2820],seed[2896],seed[2357],seed[2809],seed[3748],seed[2714],seed[3403],seed[2126],seed[2470],seed[1953],seed[2857],seed[901],seed[152],seed[3052],seed[4063],seed[3114],seed[1820],seed[3804],seed[2427],seed[2572],seed[4076],seed[1810],seed[1946],seed[2482],seed[3072],seed[1086],seed[1266],seed[1179],seed[1845],seed[479],seed[1913],seed[1085],seed[3349],seed[3955],seed[2837],seed[864],seed[2792],seed[3491],seed[705],seed[3406],seed[422],seed[3776],seed[3751],seed[456],seed[1296],seed[2555],seed[1781],seed[30],seed[3539],seed[1760],seed[2397],seed[15],seed[3790],seed[650],seed[2109],seed[929],seed[2766],seed[3143],seed[844],seed[3842],seed[2020],seed[941],seed[548],seed[3525],seed[2383],seed[911],seed[2782],seed[2901],seed[648],seed[2893],seed[620],seed[3598],seed[2543],seed[2303],seed[3896],seed[737],seed[3364],seed[3366],seed[2238],seed[1093],seed[25],seed[3159],seed[2255],seed[2327],seed[3575],seed[2159],seed[2762],seed[999],seed[3799],seed[1309],seed[1089],seed[697],seed[2356],seed[535],seed[3422],seed[528],seed[3380],seed[1990],seed[2951],seed[2731],seed[2950],seed[2877],seed[846],seed[2826],seed[843],seed[2904],seed[3750],seed[572],seed[147],seed[3822],seed[3845],seed[1515],seed[1530],seed[1524],seed[1040],seed[794],seed[2403],seed[3218],seed[3661],seed[2304],seed[3784],seed[2827],seed[3040],seed[151],seed[3151],seed[598],seed[1128],seed[748],seed[933],seed[3152],seed[499],seed[1801],seed[670],seed[3068],seed[2011],seed[776],seed[3496],seed[1730],seed[2897],seed[2274],seed[2571],seed[557],seed[1340],seed[1343],seed[2779],seed[296],seed[3623],seed[1320],seed[195],seed[3145],seed[2991],seed[3716],seed[3280],seed[3059],seed[1080],seed[2536],seed[2494],seed[730],seed[2513],seed[223],seed[443],seed[132],seed[1991],seed[2883],seed[3020],seed[1495],seed[3226],seed[1989],seed[3981],seed[1058],seed[3733],seed[2165],seed[2899],seed[3587],seed[1829],seed[4031],seed[2996],seed[584],seed[1789],seed[2056],seed[3460],seed[1498],seed[2341],seed[2040],seed[273],seed[1703],seed[3293],seed[2667],seed[625],seed[2884],seed[2852],seed[3999],seed[3540],seed[2585],seed[2359],seed[1644],seed[2484],seed[797],seed[1130],seed[2474],seed[2460],seed[3771],seed[3596],seed[3528],seed[1678],seed[3438],seed[194],seed[3638],seed[186],seed[1541],seed[565],seed[2881],seed[617],seed[531],seed[1386],seed[3829],seed[4046],seed[1082],seed[3351],seed[638],seed[820],seed[3870],seed[3046],seed[143],seed[1725],seed[372],seed[3589],seed[3936],seed[2959],seed[511],seed[1611],seed[414],seed[2353],seed[2646],seed[3416],seed[3106],seed[141],seed[4080],seed[540],seed[3212],seed[2926],seed[526],seed[1380],seed[2501],seed[3887],seed[3352],seed[3902],seed[438],seed[175],seed[2290],seed[3869],seed[1475],seed[3026],seed[809],seed[2207],seed[3608],seed[1428],seed[1956],seed[1302],seed[66],seed[189],seed[3749],seed[2451],seed[3030],seed[307],seed[2128],seed[2072],seed[2329],seed[4036],seed[2804],seed[712],seed[951],seed[3166],seed[1779],seed[3169],seed[3546],seed[1788],seed[1193],seed[3098],seed[812],seed[167],seed[2086],seed[233],seed[2479],seed[4055],seed[3696],seed[2748],seed[3332],seed[472],seed[1211],seed[4003],seed[3229],seed[1414],seed[2561],seed[2472],seed[3445],seed[2962],seed[3806],seed[1634],seed[583],seed[3242],seed[2288],seed[1571],seed[3585],seed[3358],seed[848],seed[3605],seed[524],seed[3946],seed[665],seed[3774],seed[2594],seed[3389],seed[256],seed[343],seed[509],seed[1382],seed[1529],seed[2065],seed[2395],seed[2957],seed[1777],seed[3164],seed[1695],seed[1840],seed[1148],seed[3409],seed[2085],seed[3817],seed[351],seed[1107],seed[3267],seed[788],seed[790],seed[815],seed[2314],seed[2296],seed[2631],seed[1507],seed[3126],seed[3296],seed[2887],seed[742],seed[503],seed[898],seed[3302],seed[3904],seed[60],seed[754],seed[859],seed[3300],seed[3788],seed[139],seed[1528],seed[2468],seed[3557],seed[1400],seed[1459],seed[1723],seed[3340],seed[1959],seed[1350],seed[689],seed[2704],seed[2919],seed[1387],seed[3927],seed[2999],seed[3890],seed[2993],seed[2863],seed[402],seed[3943],seed[1015],seed[2316],seed[1104],seed[169],seed[1252],seed[1714],seed[2146],seed[1011],seed[2050],seed[520],seed[3319],seed[3653],seed[2203],seed[3824],seed[408],seed[1440],seed[2791],seed[145],seed[1009],seed[1671],seed[2089],seed[106],seed[1531],seed[1006],seed[4016],seed[236],seed[1446],seed[3237],seed[2037],seed[784],seed[675],seed[914],seed[1910],seed[1969],seed[1784],seed[3787],seed[3702],seed[3093],seed[450],seed[3724],seed[3601],seed[439],seed[1927],seed[971],seed[542],seed[915],seed[1915],seed[10],seed[1154],seed[1646],seed[1743],seed[3882],seed[1463],seed[17],seed[1132],seed[943],seed[176],seed[916],seed[2564],seed[1584],seed[1883],seed[395],seed[3084],seed[3586],seed[1766],seed[1871],seed[2478],seed[107],seed[1149],seed[2133],seed[266],seed[564],seed[3550],seed[3667],seed[1171],seed[3920],seed[2839],seed[3230],seed[1720],seed[454],seed[3337],seed[2535],seed[1341],seed[1468],seed[2183],seed[2311],seed[1805],seed[3582],seed[1793],seed[1114],seed[599],seed[2438],seed[957],seed[310],seed[392],seed[3686],seed[1771],seed[3374],seed[1888],seed[3109],seed[749],seed[1493],seed[4079],seed[4017],seed[1947],seed[1162],seed[4029],seed[701],seed[82],seed[4020],seed[3011],seed[2135],seed[3997],seed[1250],seed[3618],seed[1583],seed[1694],seed[3808],seed[3819],seed[2866],seed[913],seed[397],seed[657],seed[3231],seed[821],seed[3743],seed[1467],seed[1904],seed[3958],seed[374],seed[4040],seed[3655],seed[1565],seed[3592],seed[3534],seed[3578],seed[2666],seed[2176],seed[1469],seed[3034],seed[421],seed[1259],seed[2396],seed[1778],seed[1884],seed[3669],seed[1163],seed[2394],seed[3657],seed[1677],seed[695],seed[126],seed[2261],seed[2604],seed[739],seed[1425],seed[3149],seed[2688],seed[2713],seed[2015],seed[118],seed[1988],seed[1419],seed[1828],seed[2210],seed[2652],seed[1084],seed[2355],seed[549],seed[1146],seed[2789],seed[2636],seed[740],seed[2201],seed[65],seed[1581],seed[350],seed[1216],seed[2645],seed[1851],seed[924],seed[2305],seed[2217],seed[3966],seed[4064],seed[3827],seed[1660],seed[3088],seed[2410],seed[3972],seed[1841],seed[1735],seed[587],seed[4085],seed[1473],seed[3180],seed[921],seed[2786],seed[28],seed[871],seed[1717],seed[2041],seed[3234],seed[2721],seed[434],seed[3111],seed[3041],seed[639],seed[2684],seed[3039],seed[3580],seed[1876],seed[2345],seed[644],seed[3117],seed[3531],seed[2405],seed[1023],seed[3001],seed[905],seed[3617],seed[387],seed[2254],seed[2424],seed[4073],seed[3225],seed[1487],seed[1757],seed[405],seed[3303],seed[3271],seed[3713],seed[37],seed[1397],seed[3588],seed[3726],seed[2569],seed[750],seed[1290],seed[3295],seed[2700],seed[807],seed[2680],seed[124],seed[3603],seed[1786],seed[1143],seed[359],seed[1105],seed[398],seed[340],seed[3719],seed[3100],seed[1318],seed[2349],seed[1257],seed[3912],seed[1938],seed[3915],seed[1245],seed[618],seed[2986],seed[76],seed[3547],seed[3228],seed[1905],seed[573],seed[2477],seed[3710],seed[3019],seed[681],seed[1092],seed[2491],seed[404],seed[3763],seed[1511],seed[228],seed[171],seed[727],seed[3542],seed[271],seed[677],seed[3025],seed[1638],seed[1359],seed[2368],seed[3318],seed[239],seed[746],seed[1488],seed[493],seed[3834],seed[3913],seed[708],seed[2799],seed[3768],seed[2036],seed[2229],seed[1304],seed[1534],seed[3634],seed[1598],seed[1768],seed[3988],seed[2400],seed[3621],seed[508],seed[3350],seed[2921],seed[384],seed[3077],seed[3664],seed[2755],seed[1798],seed[2105],seed[3903],seed[498],seed[658],seed[44],seed[3015],seed[3922],seed[373],seed[635],seed[1698],seed[2741],seed[1547],seed[1328],seed[1020],seed[2235],seed[1144],seed[3139],seed[2267],seed[1732],seed[324],seed[1753],seed[830],seed[1150],seed[3497],seed[39],seed[1066],seed[309],seed[2956],seed[3637],seed[487],seed[170],seed[3244],seed[3083],seed[3137],seed[3215],seed[1147],seed[481],seed[1982],seed[566],seed[2747],seed[3894],seed[2580],seed[3116],seed[1687],seed[2966],seed[2635],seed[2313],seed[1330],seed[2623],seed[462],seed[882],seed[217],seed[3720],seed[320],seed[2481],seed[1235],seed[968],seed[3256],seed[3119],seed[3830],seed[393],seed[3270],seed[731],seed[1447],seed[3888],seed[43],seed[758],seed[974],seed[2930],seed[2683],seed[483],seed[629],seed[988],seed[2240],seed[1490],seed[2891],seed[2278],seed[2697],seed[2366],seed[3835],seed[3919],seed[3604],seed[2874],seed[3217],seed[2931],seed[255],seed[2158],seed[2271],seed[806],seed[52],seed[994],seed[250],seed[1650],seed[1613],seed[3607],seed[1415],seed[1413],seed[1206],seed[2178],seed[683],seed[500],seed[3521],seed[506],seed[291],seed[3167],seed[1321],seed[2875],seed[45],seed[2964],seed[1356],seed[3078],seed[3984],seed[1029],seed[1596],seed[2450],seed[3559],seed[1748],seed[2337],seed[2272],seed[2797],seed[2344],seed[2596],seed[2695],seed[158],seed[4053],seed[1708],seed[2012],seed[3873],seed[2710],seed[2352],seed[2031],seed[2719],seed[926],seed[1228],seed[559],seed[491],seed[2894],seed[1846],seed[3619],seed[803],seed[2429],seed[1033],seed[1332],seed[3932],seed[2489],seed[1135],seed[3346],seed[2612],seed[2522],seed[2739],seed[1974],seed[1594],seed[3197],seed[3173],seed[2389],seed[1354],seed[1039],seed[856],seed[2033],seed[1960],seed[2862],seed[721],seed[3769],seed[3558],seed[2622],seed[902],seed[919],seed[3357],seed[2589],seed[153],seed[3367],seed[651],seed[3456],seed[3606],seed[959],seed[2856],seed[3459],seed[1542],seed[49],seed[4047],seed[3395],seed[4035],seed[85],seed[278],seed[1478],seed[3755],seed[168],seed[2375],seed[148],seed[369],seed[1426],seed[614],seed[245],seed[3962],seed[1633],seed[488],seed[4],seed[2581],seed[837],seed[2679],seed[2098],seed[1822],seed[347],seed[2005],seed[610],seed[3708],seed[3133],seed[981],seed[103],seed[2758],seed[1630],seed[2431],seed[3398],seed[1661],seed[3199],seed[308],seed[1286],seed[1901],seed[2851],seed[1664],seed[698],seed[1207],seed[3042],seed[2526],seed[46],seed[1849],seed[117],seed[2685],seed[1881],seed[2250],seed[3440],seed[1116],seed[3063],seed[3956],seed[1679],seed[1657],seed[3959],seed[2437],seed[1272],seed[868],seed[3208],seed[2847],seed[3421],seed[2915],seed[755],seed[2066],seed[1432],seed[2725],seed[2798],seed[218],seed[2189],seed[3467],seed[83],seed[3691],seed[3615],seed[1996],seed[3372],seed[4052],seed[2870],seed[3681],seed[3625],seed[910],seed[522],seed[3064],seed[2832],seed[1522],seed[87],seed[558],seed[702],seed[655],seed[2488],seed[411],seed[977],seed[98],seed[3986],seed[896],seed[2582],seed[474],seed[3765],seed[2780],seed[9],seed[2503],seed[3926],seed[1686],seed[162],seed[2992],seed[3251],seed[3209],seed[586],seed[2],seed[3690],seed[2273],seed[2933],seed[2961],seed[1830],seed[2074],seed[4082],seed[2726],seed[437],seed[1101],seed[976],seed[12],seed[99],seed[1158],seed[3561],seed[2563],seed[1609],seed[764],seed[105],seed[847],seed[226],seed[1295],seed[3263],seed[1247],seed[401],seed[1112],seed[964],seed[3368],seed[2480],seed[3745],seed[1159],seed[1680],seed[3954],seed[67],seed[2360],seed[2323],seed[34],seed[2161],seed[3780],seed[2293],seed[1999],seed[3150],seed[3115],seed[3742],seed[2234],seed[1872],seed[2508],seed[3654],seed[3384],seed[417],seed[406],seed[3317],seed[4050],seed[1188],seed[2407],seed[1125],seed[607],seed[2506],seed[2096],seed[950],seed[831],seed[197],seed[3732],seed[2559],seed[2978],seed[962],seed[2821],seed[3635],seed[3851],seed[2675],seed[3359],seed[3375],seed[2817],seed[79],seed[2546],seed[1591],seed[280],seed[3158],seed[2131],seed[2614],seed[2527],seed[2317],seed[1007],seed[3449],seed[2947],seed[1763],seed[2197],seed[2309],seed[3929],seed[1361],seed[747],seed[2689],seed[2960],seed[3569],seed[3016],seed[1917],seed[1852],seed[612],seed[1800],seed[711],seed[461],seed[2900],seed[383],seed[137],seed[2184],seed[2463],seed[1833],seed[1333],seed[282],seed[760],seed[3476],seed[292],seed[1357],seed[2227],seed[3644],seed[2245],seed[2315],seed[3567],seed[900],seed[3891],seed[346],seed[1976],seed[1658],seed[3797],seed[41],seed[3257],seed[3701],seed[1255],seed[1076],seed[909],seed[2139],seed[1138],seed[580],seed[1311],seed[3815],seed[3998],seed[2452],seed[1018],seed[2059],seed[1243],seed[2946],seed[1377],seed[3941],seed[1608],seed[284],seed[3793],seed[2285],seed[2208],seed[1620],seed[2114],seed[539],seed[2983],seed[2749],seed[2283],seed[3648],seed[2289],seed[925],seed[1050],seed[1293],seed[1751],seed[3683],seed[3680],seed[4004],seed[2640],seed[1482],seed[1131],seed[3849],seed[3626],seed[3233],seed[3009],seed[3189],seed[3833],seed[237],seed[116],seed[33],seed[51],seed[2542],seed[3995],seed[1503],seed[2770],seed[3005],seed[3792],seed[4008],seed[1826],seed[1886],seed[4058],seed[2340],seed[2910],seed[1019],seed[2232],seed[92],seed[330],seed[3939],seed[2935],seed[2765],seed[2505],seed[1971],seed[2660],seed[3862],seed[3832],seed[2761],seed[653],seed[3253],seed[3933],seed[3102],seed[1726],seed[341],seed[1355],seed[979],seed[2358],seed[1263],seed[619],seed[3194],seed[1706],seed[1083],seed[432],seed[1992],seed[2191],seed[2043],seed[2708],seed[2558],seed[1770],seed[453],seed[1178],seed[2544],seed[2123],seed[1450],seed[2118],seed[1232],seed[2045],seed[2231],seed[2213],seed[3854],seed[2917],seed[570],seed[21],seed[1683],seed[3688],seed[3183],seed[1065],seed[3435],seed[3415],seed[836],seed[1589],seed[2286],seed[3934],seed[1063],seed[3490],seed[3970],seed[1041],seed[814],seed[829],seed[3642],seed[932],seed[810],seed[1625],seed[792],seed[1607],seed[3004],seed[1891],seed[2672],seed[2302],seed[756],seed[1755],seed[2029],seed[3043],seed[2369],seed[736],seed[4056],seed[1604],seed[2433],seed[1847],seed[2705],seed[2734],seed[270],seed[3092],seed[2912],seed[283],seed[3612],seed[1856],seed[2476],seed[2858],seed[2785],seed[3283],seed[2663],seed[2905],seed[1616],seed[2590],seed[3455],seed[2702],seed[3419],seed[2025],seed[884],seed[3472],seed[1574],seed[1642],seed[533],seed[2754],seed[3014],seed[2764],seed[543],seed[2225],seed[728],seed[2583],seed[879],seed[2101],seed[1021],seed[1168],seed[918],seed[3649],seed[538],seed[1564],seed[1056],seed[1759],seed[1705],seed[4092],seed[1456],seed[3568],seed[2143],seed[3205],seed[2462],seed[2243],seed[2613],seed[2370],seed[707],seed[2443],seed[1170],seed[1980],seed[779],seed[135],seed[2063],seed[1544],seed[187],seed[3241],seed[3436],seed[2046],seed[2952],seed[3679],seed[3177],seed[2658],seed[262],seed[1003],seed[1268],seed[1152],seed[2330],seed[2639],seed[2198],seed[2413],seed[1662],seed[1472],seed[1395],seed[164],seed[1807],seed[823],seed[2846],seed[3309],seed[96],seed[2321],seed[723],seed[673],seed[2090],seed[716],seed[656],seed[2144],seed[2694],seed[1769],seed[2112],seed[1283],seed[1237],seed[3731],seed[2554],seed[3982],seed[2385],seed[1920],seed[832],seed[1525],seed[956],seed[636],seed[4091],seed[285],seed[3447],seed[1555],seed[1970],seed[1639],seed[936],seed[2822],seed[1823],seed[1265],seed[609],seed[1827],seed[1692],seed[3345],seed[2172],seed[337],seed[3272],seed[1615],seed[1612],seed[3508],seed[3899],seed[2584],seed[2038],seed[883],seed[3338],seed[1722],seed[3573],seed[996],seed[3138],seed[1587],seed[322],seed[3101],seed[972],seed[2932],seed[3124],seed[1127],seed[91],seed[1017],seed[726],seed[3944],seed[459],seed[2953],seed[628],seed[1814],seed[2740],seed[2001],seed[3344],seed[2148],seed[2654],seed[3067],seed[281],seed[2265],seed[2752],seed[778],seed[3090],seed[2855],seed[2416],seed[3636],seed[1684],seed[863],seed[269],seed[1307],seed[3965],seed[3390],seed[3747],seed[3323],seed[2391],seed[3376],seed[1973],seed[198],seed[2840],seed[3045],seed[2280],seed[3182],seed[2968],seed[2763],seed[983],seed[1649],seed[2019],seed[265],seed[3548],seed[1059],seed[1669],seed[3712],seed[1067],seed[3831],seed[1838],seed[2399],seed[2609],seed[3692],seed[2818],seed[3154],seed[1517],seed[2669],seed[354],seed[3689],seed[3356],seed[389],seed[1399],seed[1457],seed[1572],seed[2387],seed[3037],seed[1621],seed[2174],seed[2498],seed[2963],seed[2872],seed[2574],seed[3495],seed[1433],seed[3898],seed[1546],seed[2934],seed[2469],seed[2032],seed[1809],seed[2196],seed[992],seed[3600],seed[514],seed[714],seed[183],seed[2325],seed[3107],seed[3140],seed[3450],seed[111],seed[771],seed[920],seed[1254],seed[2743],seed[3289],seed[970],seed[3299],seed[3990],seed[2618],seed[3171],seed[3878],seed[3532],seed[2129],seed[1052],seed[3439],seed[1889],seed[889],seed[504],seed[2119],seed[364],seed[1367],seed[306],seed[3584],seed[3204],seed[4054],seed[822],seed[370],seed[3314],seed[1212],seed[2435],seed[2751],seed[3168],seed[2716],seed[1729],seed[1986],seed[2729],seed[3315],seed[3412],seed[261],seed[3857],seed[1069],seed[4078],seed[547],seed[3816],seed[1198],seed[2655],seed[3994],seed[3960],seed[1995],seed[2047],seed[1958],seed[295],seed[4012],seed[3091],seed[3400],seed[1000],seed[264],seed[1427],seed[1124],seed[562],seed[3501],seed[594],seed[1203],seed[1253],seed[2116],seed[2637],seed[154],seed[980],seed[2257],seed[1412],seed[3482],seed[3473],seed[732],seed[3694],seed[2153],seed[1627],seed[2674],seed[1269],seed[2351],seed[1389],seed[2166],seed[1392],seed[3576],seed[2981],seed[4039],seed[352],seed[2262],seed[3477],seed[26],seed[2511],seed[1962],seed[3062],seed[316],seed[3825],seed[2336],seed[1274],seed[1641],seed[1194],seed[215],seed[2379],seed[2647],seed[3393],seed[3408],seed[144],seed[3511],seed[2287],seed[1563],seed[928],seed[3122],seed[1273],seed[3307],seed[62],seed[3500],seed[201],seed[1911],seed[2319],seed[2732],seed[2718],seed[1939],seed[1081],seed[2914],seed[1480],seed[3821],seed[214],seed[1853],seed[3335],seed[2744],seed[1022],seed[2458],seed[1994],seed[3292],seed[3783],seed[3807],seed[2717],seed[4088],seed[104],seed[3488],seed[3693],seed[912],seed[2682],seed[4000],seed[263],seed[1032],seed[1176],seed[2595],seed[874],seed[3021],seed[2414],seed[1984],seed[780],seed[2099],seed[632],seed[138],seed[3761],seed[3530],seed[2568],seed[569],seed[2841],seed[1998],seed[3852],seed[2879],seed[3287],seed[1455],seed[1737],seed[3746],seed[3897],seed[2266],seed[2211],seed[14],seed[1102],seed[334],seed[2268],seed[1783],seed[507],seed[2607],seed[3252],seed[3803],seed[1854],seed[363],seed[2392],seed[3647],seed[1383],seed[2845],seed[1817],seed[3076],seed[379],seed[2529],seed[478],seed[1552],seed[19],seed[3916],seed[1665],seed[1600],seed[1445],seed[1349],seed[1700],seed[2814],seed[2989],seed[1486],seed[3007],seed[3110],seed[965],seed[2892],seed[323],seed[3254],seed[1937],seed[800],seed[1504],seed[4014],seed[3103],seed[603],seed[1120],seed[907],seed[2880],seed[1197],seed[2256],seed[1610],seed[944],seed[2120],seed[179],seed[3483],seed[1028],seed[4032],seed[1727],seed[3554],seed[1746],seed[3938],seed[942],seed[1586],seed[234],seed[1559],seed[2500],seed[2578],seed[484],seed[2771],seed[3715],seed[3160],seed[1371],seed[3855],seed[3651],seed[3505],seed[3645],seed[1844],seed[2502],seed[1261],seed[2298],seed[530],seed[3373],seed[2269],seed[74],seed[333],seed[3250],seed[1954],seed[3678],seed[1799],seed[2067],seed[3658],seed[849],seed[2911],seed[1711],seed[3814],seed[3652],seed[394],seed[3261],seed[3973],seed[1270],seed[1164],seed[3992],seed[1182],seed[3097],seed[205],seed[2677],seed[2170],seed[3249],seed[140],seed[428],seed[3969],seed[3430],seed[1606],seed[110],seed[1064],seed[409],seed[3730],seed[2062],seed[2634],seed[2854],seed[947],seed[299],seed[114],seed[1520],seed[182],seed[2998],seed[3222],seed[2549],seed[246],seed[329],seed[3650],seed[3207],seed[3509],seed[2324],seed[1209],seed[2520],seed[1481],seed[2361],seed[275],seed[2057],seed[2013],seed[468],seed[1190],seed[1129],seed[1411],seed[1260],seed[568],seed[2530],seed[2111],seed[1294],seed[687],seed[469],seed[1957],seed[431],seed[2515],seed[1819],seed[691],seed[3232],seed[3964],seed[880],seed[2601],seed[178],seed[3434],seed[1908],seed[786],seed[2657],seed[805],seed[2068],seed[2617],seed[1218],seed[3820],seed[2805],seed[4026],seed[1460],seed[1204],seed[1435],seed[1024],seed[2728],seed[3413],seed[2916],seed[2204],seed[3392],seed[2838],seed[181],seed[2404],seed[1929],seed[2200],seed[1313],seed[3562],seed[1142],seed[1483],seed[423],seed[3924],seed[3443],seed[1690],seed[1035],seed[505],seed[2816],seed[2665],seed[774],seed[4049],seed[2735],seed[2547],seed[1569],seed[1443],seed[2382],seed[984],seed[1987],seed[88],seed[1244],seed[841],seed[987],seed[3759],seed[358],seed[1774],seed[1602],seed[525],seed[2597],seed[400],seed[4048],seed[2643],seed[3262],seed[704],seed[3752],seed[674],seed[2775],seed[1979],seed[1935],seed[2651],seed[3910],seed[3288],seed[2260],seed[3044],seed[516],seed[35],seed[2007],seed[150],seed[1985],seed[855],seed[3739],seed[862],seed[2670],seed[2457],seed[3850],seed[903],seed[1477],seed[3074],seed[789],seed[327],seed[2727],seed[1636],seed[3671],seed[311],seed[1369],seed[3672],seed[3662],seed[78],seed[2599],seed[3094],seed[873],seed[2556],seed[2737],seed[2552],seed[3753],seed[1496],seed[3457],seed[2707],seed[3125],seed[1754],seed[1298],seed[1351],seed[317],seed[466],seed[3027],seed[3087],seed[2378],seed[1097],seed[3949],seed[1739],seed[1335],seed[1526],seed[3876],seed[2698],seed[1401],seed[3404],seed[1205],seed[2514],seed[3564],seed[899],seed[480],seed[209],seed[4090],seed[1712],seed[3828],seed[678],seed[2955],seed[1718],seed[2690],seed[1704],seed[865],seed[1601],seed[2028],seed[3722],seed[2440],seed[1462],seed[3754],seed[2807],seed[3853],seed[3070],seed[2372],seed[767],seed[2709],seed[1812],seed[3794],seed[2426],seed[1217],seed[2276],seed[2860],seed[3475],seed[2678],seed[1775],seed[1342],seed[3035],seed[2850],seed[2490],seed[2745],seed[2363],seed[2475],seed[1436],seed[1652],seed[3581],seed[3361],seed[3095],seed[819],seed[3360],seed[2228],seed[2746],seed[1925],seed[3487],seed[303],seed[1590],seed[1691],seed[3844],seed[1707],seed[2455],seed[1635],seed[2813],seed[791],seed[180],seed[934],seed[1818],seed[2808],seed[2075],seed[2083],seed[272],seed[2155],seed[1037],seed[452],seed[2466],seed[289],seed[3555],seed[751],seed[2519],seed[294],seed[606],seed[3130],seed[3494],seed[2423],seed[2898],seed[709],seed[349],seed[2122],seed[120],seed[3484],seed[4093],seed[3146],seed[816],seed[3333],seed[3577],seed[2331],seed[2456],seed[1562],seed[3128],seed[3071],seed[1258],seed[738],seed[61],seed[649],seed[2308],seed[216],seed[1416],seed[4019],seed[923],seed[1157],seed[1899],seed[3885],seed[2149],seed[3216],seed[998],seed[3989],seed[3336],seed[3433],seed[319],seed[2027],seed[1264],seed[68],seed[1281],seed[672],seed[1685],seed[596],seed[799],seed[326],seed[1249],seed[3474],seed[161],seed[2975],seed[3310],seed[930],seed[2428],seed[3381],seed[940],seed[866],seed[510],seed[3524],seed[3414],seed[2493],seed[2800],seed[3134],seed[3823],seed[2611],seed[1967],seed[3945],seed[24],seed[2087],seed[2687],seed[954],seed[1016],seed[3423],seed[2365],seed[3000],seed[2742],seed[1936],seed[1997],seed[637],seed[1538],seed[3008],seed[3179],seed[2783],seed[3940],seed[1471],seed[3112],seed[1172],seed[1417],seed[1223],seed[2539],seed[3326],seed[3363],seed[3613],seed[604],seed[2364],seed[1628],seed[3947],seed[818],seed[613],seed[4028],seed[3796],seed[1444],seed[2377],seed[3113],seed[1381],seed[3266],seed[206],seed[1857],seed[783],seed[3033],seed[2186],seed[3424],seed[4062],seed[1238],seed[512],seed[1122],seed[5],seed[220],seed[1902],seed[1167],seed[2081],seed[84],seed[1894],seed[22],seed[494],seed[1756],seed[4001],seed[1113],seed[3468],seed[2060],seed[2134],seed[2249],seed[2000],seed[2284],seed[2824],seed[2140],seed[1378],seed[948],seed[3843],seed[1548],seed[3135],seed[1580],seed[1213],seed[1912],seed[1792],seed[251],seed[3198],seed[2064],seed[840],seed[2002],seed[2310],seed[1345],seed[845],seed[534],seed[2322],seed[2843],seed[2889],seed[1096],seed[995],seed[2603],seed[2194],seed[1161],seed[254],seed[298],seed[4030],seed[1697],seed[3486],seed[3089],seed[2819],seed[55],seed[377],seed[2496],seed[3781],seed[1236],seed[260],seed[1681],seed[890],seed[2938],seed[3418],seed[36],seed[32],seed[3304],seed[1539],seed[1568],seed[1241],seed[360],seed[2659],seed[1423],seed[2242],seed[1922],seed[743],seed[2936],seed[2039],seed[3493],seed[2082],seed[682],seed[3297],seed[1721],seed[757],seed[1592],seed[3921],seed[2388],seed[314],seed[3925],seed[2073],seed[290],seed[2518],seed[852],seed[2320],seed[3277],seed[3991],seed[227],seed[1532],seed[396],seed[258],seed[1859],seed[2965],seed[949],seed[2925],seed[1951],seed[2292],seed[1422],seed[2949],seed[3627],seed[366],seed[1476],seed[447],seed[1710],seed[1863],seed[601],seed[661],seed[3099],seed[1347],seed[1300],seed[1322],seed[3778],seed[2010],seed[3017],seed[1808],seed[835],seed[1848],seed[627],seed[1312],seed[1659],seed[2248],seed[667],seed[3536],seed[1667],seed[27],seed[2873],seed[2104],seed[766],seed[2448],seed[654],seed[2219],seed[2830],seed[355],seed[1752],seed[448],seed[2160],seed[365],seed[3196],seed[1325],seed[706],seed[3331],seed[427],seed[3362],seed[1156],seed[1110],seed[1868],seed[3162],seed[2202],seed[3704],seed[121],seed[1963],seed[2650],seed[1437],seed[3471],seed[3616],seed[4057],seed[2053],seed[1474],seed[3723],seed[1595],seed[3928],seed[399],seed[2630],seed[3085],seed[2142],seed[1787],seed[3838],seed[3282],seed[722],seed[878],seed[1222],seed[3677],seed[1484],seed[3812],seed[149],seed[3224],seed[1764],seed[1508],seed[2220],seed[2301],seed[616],seed[204],seed[119],seed[2693],seed[1839],seed[1470],seed[1410],seed[2902],seed[2354],seed[734],seed[1897],seed[1215],seed[735],seed[3161],seed[230],seed[3328],seed[2720],seed[666],seed[860],seed[2886],seed[1513],seed[3560],seed[2077],seed[2214],seed[185],seed[985],seed[58],seed[3239],seed[305],seed[3410],seed[1825],seed[3777],seed[1981],seed[3308],seed[1174],seed[1358],seed[3458],seed[3245],seed[1242],seed[546],seed[2773],seed[3685],seed[2106],seed[3673],seed[477],seed[2137],seed[446],seed[1137],seed[1119],seed[3633],seed[3985],seed[416],seed[2026],seed[163],seed[893],seed[3979],seed[2927],seed[2224],seed[3371],seed[2156],seed[1299],seed[412],seed[208],seed[102],seed[2533],seed[2924],seed[1952],seed[3758],seed[2124],seed[3744],seed[1588],seed[1],seed[336],seed[2869],seed[3255],seed[2439],seed[2828],seed[1336],seed[221],seed[3656],seed[3061],seed[495],seed[2523],seed[1087],seed[3837],seed[1918],seed[2633],seed[224],seed[1219],seed[2795],seed[3451],seed[2417],seed[692],seed[2920],seed[3334],seed[3798],seed[1166],seed[3023],seed[660],seed[602],seed[1060],seed[811],seed[1944],seed[1579],seed[1452],seed[2147],seed[2509],seed[527],seed[2328],seed[4005],seed[1277],seed[643],seed[1071],seed[2668],seed[332],seed[2738],seed[2069],seed[1090],seed[3185],seed[257],seed[1797],seed[1734],seed[1696],seed[1914],seed[1656],seed[2586],seed[1407],seed[645],seed[1115],seed[1047],seed[2246],seed[1724],seed[1103],seed[2023],seed[3060],seed[579],seed[1136],seed[2138],seed[2006],seed[1536],seed[908],seed[2239],seed[1062],seed[3968],seed[4024],seed[2408],seed[94],seed[857],seed[541],seed[588],seed[2541],seed[441],seed[3327],seed[710],seed[2335],seed[1306],seed[3923],seed[1898],seed[86],seed[3846],seed[2182],seed[2548],seed[1834],seed[1108],seed[442],seed[418],seed[1314],seed[2768],seed[501],seed[2835],seed[1271],seed[2810],seed[3273],seed[2793],seed[3883],seed[664],seed[2190],seed[3847],seed[356],seed[1749],seed[241],seed[2985],seed[1034],seed[2723],seed[2163],seed[3142],seed[824],seed[939],seed[2895],seed[2421],seed[3489],seed[1042],seed[3243],seed[277],seed[3190],seed[1934],seed[2049],seed[3051],seed[3670],seed[3013],seed[3556],seed[825],seed[798],seed[1200],seed[2071],seed[3565],seed[715],seed[2903],seed[891],seed[4007],seed[1835],seed[242],seed[338],seed[3503],seed[3737],seed[93],seed[1738],seed[4089],seed[1500],seed[621],seed[1492],seed[3417],seed[2409],seed[1373],seed[2712],seed[2487],seed[1648],seed[267],seed[1663],seed[3246],seed[1645],seed[2374],seed[1765],seed[935],seed[2164],seed[4069],seed[3772],seed[3735],seed[403],seed[225],seed[1877],seed[4023],seed[13],seed[1892],seed[3782],seed[3105],seed[3545],seed[3341],seed[4068],seed[1831],seed[2878],seed[3452],seed[3120],seed[1118],seed[1348],seed[1326],seed[2971],seed[2467],seed[3533],seed[1449],seed[81],seed[615],seed[3498],seed[1285],seed[391],seed[3665],seed[3276],seed[3516],seed[2802],seed[3170],seed[279],seed[741],seed[3428],seed[2177],seed[1282],seed[3909],seed[3055],seed[440],seed[817],seed[1668],seed[1431],seed[2212],seed[4044],seed[293],seed[3886],seed[556],seed[1424],seed[3628],seed[2411],seed[2373],seed[4071],seed[2030],seed[1374],seed[1331],seed[2567],seed[232],seed[3200],seed[986],seed[2209],seed[57],seed[626],seed[3394],seed[519],seed[2434],seed[2620],seed[1943],seed[449],seed[759],seed[2042],seed[2598],seed[157],seed[630],seed[1715],seed[3911],seed[1699],seed[174],seed[1141],seed[1079],seed[3446],seed[1619],seed[3108],seed[2384],seed[75],seed[2094],seed[70],seed[2778],seed[1191],seed[978],seed[3227],seed[2270],seed[2815],seed[3900],seed[1790],seed[2222],seed[2662],seed[3248],seed[3721],seed[4042],seed[3397],seed[2653],seed[3339],seed[3593],seed[576],seed[128],seed[2236],seed[2141],seed[696],seed[567],seed[3786],seed[1391],seed[917],seed[435],seed[313],seed[724],seed[1094],seed[1545],seed[1945],seed[1966],seed[1240],seed[1843],seed[1933],seed[3235],seed[3330],seed[1975],seed[3544],seed[2393],seed[335],seed[1453],seed[1728],seed[3301],seed[3313],seed[1173],seed[2656],seed[3957],seed[2430],seed[1570],seed[2022],seed[3024],seed[1117],seed[2247],seed[2759],seed[1497],seed[3879],seed[1855],seed[115],seed[430],seed[1078],seed[3206],seed[966],seed[3080],seed[894],seed[1585],seed[690],seed[1519],seed[518],seed[1575],seed[1556],seed[1346],seed[1214],seed[4061],seed[600],seed[4083],seed[2772],seed[2722],seed[3155],seed[424],seed[3407],seed[2638],seed[318],seed[938],seed[231],seed[781],seed[1139],seed[4009],seed[3700],seed[2540],seed[961],seed[1509],seed[3574],seed[382],seed[3520],seed[173],seed[297],seed[2483],seed[2230],seed[1192],seed[3874],seed[1398],seed[719],seed[3538],seed[1091],seed[1907],seed[1100],seed[2787],seed[3875],seed[2088],seed[2079],seed[858],seed[3469],seed[2115],seed[253],seed[536],seed[1861],seed[1761],seed[1442],seed[3279],seed[2908],seed[881],seed[3948],seed[3935],seed[2608],seed[3213],seed[3795],seed[3741],seed[3674],seed[2550],seed[3427],seed[1647],seed[2923],seed[4094],seed[429],seed[1670],seed[1491],seed[1896],seed[1439],seed[993],seed[1368],seed[2241],seed[1388],seed[2497],seed[445],seed[1464],seed[3465],seed[2127],seed[1693],seed[1521],seed[853],seed[3184],seed[2080],seed[2906],seed[11],seed[3378],seed[1134],seed[2048],seed[2380],seed[134],seed[3385],seed[2984],seed[1025],seed[1220],seed[4018],seed[3066],seed[2537],seed[1502],seed[1195]}),
        .cross_prob(cross_prob),
        .codeword(codeword10),
        .received(received10)
        );
    
    bsc bsc11(
        .clk(clk),
        .reset(reset),
        .seed({seed[3087],seed[1951],seed[3590],seed[2376],seed[2635],seed[2218],seed[1822],seed[1923],seed[2732],seed[2860],seed[4086],seed[1029],seed[797],seed[1074],seed[2774],seed[2625],seed[338],seed[240],seed[616],seed[1283],seed[2368],seed[3039],seed[2562],seed[2865],seed[3375],seed[3057],seed[1999],seed[2116],seed[2823],seed[907],seed[856],seed[3847],seed[1514],seed[535],seed[1625],seed[2983],seed[807],seed[2746],seed[2113],seed[2094],seed[2434],seed[25],seed[1781],seed[2951],seed[1607],seed[1349],seed[1420],seed[3242],seed[3770],seed[2520],seed[1593],seed[1931],seed[1520],seed[1597],seed[3310],seed[1161],seed[813],seed[1571],seed[1254],seed[172],seed[3474],seed[2550],seed[609],seed[677],seed[2314],seed[2490],seed[3977],seed[1736],seed[3223],seed[2748],seed[1783],seed[1044],seed[2229],seed[3060],seed[3093],seed[2590],seed[3976],seed[1078],seed[1009],seed[2345],seed[1744],seed[1899],seed[2986],seed[2799],seed[660],seed[2680],seed[1488],seed[3448],seed[1250],seed[2270],seed[2644],seed[2928],seed[2016],seed[1582],seed[2864],seed[744],seed[2688],seed[66],seed[435],seed[2427],seed[2243],seed[2197],seed[1090],seed[720],seed[546],seed[689],seed[1057],seed[2668],seed[3490],seed[143],seed[2265],seed[2672],seed[2831],seed[2227],seed[2977],seed[1836],seed[1286],seed[270],seed[2666],seed[3081],seed[93],seed[1769],seed[3903],seed[787],seed[668],seed[1140],seed[750],seed[2948],seed[1155],seed[3211],seed[1208],seed[1831],seed[1542],seed[3673],seed[2740],seed[1144],seed[1911],seed[1847],seed[2246],seed[3067],seed[2226],seed[937],seed[190],seed[2964],seed[1894],seed[2463],seed[3182],seed[2884],seed[3792],seed[1401],seed[3311],seed[2881],seed[3410],seed[2543],seed[1060],seed[1065],seed[1468],seed[2082],seed[3188],seed[2849],seed[2322],seed[2030],seed[2443],seed[1082],seed[2420],seed[656],seed[265],seed[669],seed[685],seed[3080],seed[3281],seed[1369],seed[3734],seed[1383],seed[3010],seed[786],seed[3822],seed[636],seed[706],seed[3716],seed[132],seed[289],seed[2652],seed[1404],seed[2608],seed[1709],seed[3818],seed[1915],seed[432],seed[1100],seed[1224],seed[3777],seed[1813],seed[1338],seed[3220],seed[3917],seed[323],seed[2177],seed[2988],seed[2425],seed[247],seed[3268],seed[3398],seed[2313],seed[3863],seed[271],seed[124],seed[931],seed[1367],seed[2927],seed[3336],seed[407],seed[3459],seed[1977],seed[1213],seed[3186],seed[1305],seed[1067],seed[3204],seed[2115],seed[593],seed[3196],seed[2004],seed[1463],seed[2843],seed[3497],seed[3425],seed[1527],seed[905],seed[1710],seed[173],seed[2727],seed[1106],seed[2891],seed[2650],seed[2255],seed[3820],seed[3450],seed[3812],seed[625],seed[885],seed[1869],seed[2319],seed[2236],seed[886],seed[2228],seed[3793],seed[419],seed[1059],seed[178],seed[2930],seed[1551],seed[1395],seed[1350],seed[754],seed[2579],seed[1154],seed[3114],seed[2708],seed[1688],seed[153],seed[439],seed[3833],seed[3896],seed[2918],seed[1947],seed[1695],seed[332],seed[3250],seed[315],seed[1393],seed[3680],seed[1623],seed[2366],seed[1902],seed[2971],seed[2118],seed[2885],seed[3807],seed[2158],seed[48],seed[1874],seed[680],seed[227],seed[694],seed[84],seed[3049],seed[2714],seed[3688],seed[2687],seed[881],seed[3419],seed[3249],seed[3408],seed[200],seed[4014],seed[2200],seed[2621],seed[958],seed[16],seed[1330],seed[1039],seed[1760],seed[2237],seed[3644],seed[1403],seed[3523],seed[2061],seed[1515],seed[3699],seed[3533],seed[3502],seed[945],seed[2767],seed[3938],seed[2258],seed[1197],seed[2710],seed[3888],seed[1052],seed[857],seed[1231],seed[957],seed[3981],seed[2433],seed[1870],seed[1741],seed[2093],seed[2282],seed[1457],seed[3422],seed[619],seed[101],seed[0],seed[1794],seed[3233],seed[1578],seed[507],seed[1660],seed[3526],seed[1761],seed[882],seed[3573],seed[443],seed[3035],seed[2069],seed[236],seed[1469],seed[329],seed[168],seed[421],seed[1739],seed[1963],seed[1969],seed[1236],seed[3693],seed[1091],seed[3064],seed[301],seed[2701],seed[3548],seed[2691],seed[798],seed[2402],seed[2707],seed[3234],seed[2508],seed[3996],seed[513],seed[2762],seed[2492],seed[3254],seed[3559],seed[738],seed[3287],seed[2190],seed[243],seed[1827],seed[2365],seed[1173],seed[1156],seed[2855],seed[3151],seed[2092],seed[1503],seed[588],seed[1748],seed[2169],seed[2527],seed[2330],seed[461],seed[1323],seed[503],seed[1712],seed[3909],seed[1244],seed[1331],seed[2664],seed[2578],seed[836],seed[1717],seed[1664],seed[3300],seed[3374],seed[2699],seed[1662],seed[912],seed[2803],seed[3098],seed[3338],seed[795],seed[2337],seed[2937],seed[3185],seed[2396],seed[721],seed[534],seed[948],seed[708],seed[3252],seed[3208],seed[2347],seed[2769],seed[2292],seed[2859],seed[1716],seed[76],seed[966],seed[2238],seed[2995],seed[875],seed[2819],seed[2346],seed[1816],seed[1587],seed[2468],seed[2239],seed[701],seed[2060],seed[1924],seed[2012],seed[2528],seed[3030],seed[2360],seed[1158],seed[1215],seed[1528],seed[3457],seed[2309],seed[207],seed[3293],seed[3381],seed[2730],seed[3210],seed[972],seed[141],seed[3574],seed[434],seed[3106],seed[541],seed[1055],seed[3779],seed[3462],seed[3823],seed[922],seed[1363],seed[2567],seed[1177],seed[2340],seed[437],seed[41],seed[1989],seed[902],seed[691],seed[2025],seed[3386],seed[2268],seed[455],seed[2382],seed[2580],seed[2168],seed[1202],seed[206],seed[898],seed[108],seed[852],seed[1324],seed[3889],seed[1719],seed[194],seed[2195],seed[3238],seed[2599],seed[3536],seed[122],seed[1497],seed[3356],seed[2614],seed[2934],seed[3253],seed[2047],seed[2291],seed[220],seed[2601],seed[4030],seed[1512],seed[4059],seed[2645],seed[5],seed[1807],seed[2775],seed[3984],seed[3277],seed[2872],seed[3218],seed[468],seed[1507],seed[3148],seed[341],seed[2355],seed[1178],seed[2682],seed[1088],seed[878],seed[3668],seed[1408],seed[2096],seed[2690],seed[2628],seed[3513],seed[1934],seed[3146],seed[2811],seed[2956],seed[1269],seed[1170],seed[1801],seed[1113],seed[2377],seed[1960],seed[3529],seed[3470],seed[1336],seed[1282],seed[3487],seed[556],seed[3028],seed[831],seed[695],seed[1653],seed[648],seed[217],seed[3610],seed[2828],seed[43],seed[339],seed[768],seed[3364],seed[1583],seed[2479],seed[2585],seed[3525],seed[3906],seed[318],seed[1255],seed[3550],seed[3138],seed[26],seed[2077],seed[2009],seed[1412],seed[3388],seed[2893],seed[3316],seed[2801],seed[2406],seed[2835],seed[523],seed[2968],seed[3508],seed[2279],seed[2572],seed[1204],seed[2136],seed[1610],seed[1038],seed[3290],seed[994],seed[1217],seed[3510],seed[3436],seed[1428],seed[911],seed[3011],seed[2633],seed[3911],seed[3446],seed[2328],seed[1212],seed[1049],seed[1141],seed[1838],seed[3702],seed[3578],seed[3475],seed[2686],seed[4068],seed[1810],seed[110],seed[1536],seed[3382],seed[568],seed[2189],seed[1697],seed[2401],seed[2233],seed[2250],seed[672],seed[1480],seed[3163],seed[1313],seed[1658],seed[1157],seed[3541],seed[801],seed[575],seed[4026],seed[2700],seed[773],seed[557],seed[973],seed[377],seed[1132],seed[397],seed[819],seed[4043],seed[1203],seed[2208],seed[2657],seed[1600],seed[3484],seed[1419],seed[152],seed[245],seed[3278],seed[2674],seed[2491],seed[2219],seed[2153],seed[55],seed[1601],seed[3391],seed[3222],seed[3625],seed[2648],seed[2742],seed[3308],seed[2834],seed[412],seed[3275],seed[3582],seed[3442],seed[1855],seed[3692],seed[3885],seed[1133],seed[743],seed[1853],seed[942],seed[3133],seed[3841],seed[2901],seed[1438],seed[3379],seed[3845],seed[2825],seed[29],seed[848],seed[3443],seed[2619],seed[2387],seed[1421],seed[1517],seed[510],seed[3890],seed[325],seed[985],seed[2119],seed[3628],seed[1817],seed[1056],seed[1168],seed[2217],seed[3344],seed[330],seed[46],seed[757],seed[401],seed[1939],seed[2157],seed[361],seed[1406],seed[1701],seed[1698],seed[2424],seed[4007],seed[698],seed[3198],seed[4058],seed[3961],seed[1198],seed[2352],seed[3922],seed[3272],seed[3972],seed[1543],seed[1700],seed[3165],seed[3875],seed[2139],seed[969],seed[3740],seed[2059],seed[2594],seed[1477],seed[3848],seed[1071],seed[1627],seed[4063],seed[2498],seed[1879],seed[3763],seed[1998],seed[2669],seed[1342],seed[1117],seed[2416],seed[250],seed[2461],seed[293],seed[3018],seed[3866],seed[1092],seed[2404],seed[3825],seed[1859],seed[224],seed[612],seed[747],seed[4018],seed[335],seed[1549],seed[1928],seed[1353],seed[3140],seed[3147],seed[884],seed[2904],seed[3775],seed[4047],seed[149],seed[452],seed[2781],seed[1301],seed[2362],seed[1704],seed[3506],seed[3321],seed[1464],seed[955],seed[967],seed[3879],seed[2902],seed[3636],seed[2123],seed[1222],seed[4019],seed[1162],seed[3561],seed[2386],seed[1667],seed[1793],seed[3608],seed[1680],seed[3413],seed[2180],seed[1247],seed[133],seed[587],seed[1945],seed[13],seed[2676],seed[2571],seed[2028],seed[815],seed[2378],seed[2138],seed[1315],seed[3320],seed[1965],seed[765],seed[2761],seed[3751],seed[904],seed[1436],seed[1973],seed[1297],seed[779],seed[1192],seed[258],seed[482],seed[2288],seed[628],seed[2205],seed[2895],seed[1278],seed[1196],seed[3135],seed[1509],seed[286],seed[563],seed[3919],seed[1252],seed[1656],seed[1304],seed[1339],seed[59],seed[3167],seed[756],seed[1502],seed[572],seed[722],seed[2379],seed[1239],seed[3373],seed[2867],seed[2494],seed[1575],seed[1399],seed[2369],seed[2220],seed[724],seed[1312],seed[1351],seed[3784],seed[2080],seed[538],seed[3161],seed[1833],seed[3748],seed[1111],seed[209],seed[2310],seed[2040],seed[3685],seed[3362],seed[488],seed[2500],seed[2182],seed[1755],seed[959],seed[2400],seed[1063],seed[415],seed[2752],seed[1628],seed[204],seed[3988],seed[591],seed[3819],seed[2763],seed[2114],seed[2445],seed[2336],seed[1216],seed[3332],seed[2624],seed[1424],seed[203],seed[371],seed[1279],seed[3665],seed[639],seed[3267],seed[1040],seed[277],seed[3957],seed[617],seed[1830],seed[2364],seed[1839],seed[4006],seed[2496],seed[1579],seed[3766],seed[2058],seed[979],seed[1182],seed[1249],seed[2531],seed[1335],seed[3318],seed[2980],seed[4055],seed[584],seed[1572],seed[3724],seed[2050],seed[2423],seed[1577],seed[3342],seed[3966],seed[4090],seed[3058],seed[2470],seed[2792],seed[734],seed[991],seed[2514],seed[586],seed[296],seed[2609],seed[3444],seed[2501],seed[1584],seed[1455],seed[2861],seed[3472],seed[2512],seed[350],seed[2539],seed[2641],seed[1373],seed[1861],seed[3681],seed[1083],seed[3645],seed[242],seed[3224],seed[3517],seed[2517],seed[1409],seed[281],seed[1491],seed[3024],seed[462],seed[2341],seed[1532],seed[2737],seed[1261],seed[3677],seed[626],seed[2043],seed[279],seed[1670],seed[3746],seed[1445],seed[543],seed[3191],seed[316],seed[1745],seed[598],seed[3756],seed[1073],seed[2909],seed[1903],seed[1325],seed[3121],seed[2804],seed[2758],seed[897],seed[302],seed[1955],seed[1362],seed[599],seed[3285],seed[15],seed[3447],seed[3619],seed[2155],seed[2034],seed[3044],seed[1019],seed[19],seed[3799],seed[771],seed[72],seed[1030],seed[1461],seed[566],seed[3393],seed[2171],seed[3893],seed[2906],seed[2681],seed[1268],seed[4085],seed[3181],seed[2485],seed[38],seed[2176],seed[1416],seed[3117],seed[711],seed[3205],seed[3542],seed[3059],seed[2592],seed[1322],seed[2962],seed[365],seed[1865],seed[1636],seed[1620],seed[2894],seed[3498],seed[1103],seed[60],seed[2754],seed[3209],seed[1237],seed[478],seed[2502],seed[3183],seed[1129],seed[3515],seed[363],seed[3620],seed[870],seed[3461],seed[1518],seed[1771],seed[638],seed[3778],seed[3020],seed[1715],seed[834],seed[2163],seed[3760],seed[3296],seed[675],seed[3733],seed[950],seed[2534],seed[2837],seed[2407],seed[2221],seed[8],seed[3331],seed[3309],seed[3108],seed[2278],seed[1242],seed[627],seed[3495],seed[1529],seed[849],seed[3325],seed[3654],seed[3271],seed[4020],seed[2982],seed[1631],seed[1863],seed[2194],seed[1886],seed[3789],seed[1702],seed[233],seed[3232],seed[1824],seed[2390],seed[1589],seed[883],seed[1504],seed[1022],seed[491],seed[234],seed[2908],seed[2515],seed[3759],seed[2342],seed[2991],seed[2356],seed[2032],seed[2544],seed[1691],seed[1214],seed[3951],seed[2844],seed[3174],seed[2324],seed[1265],seed[3967],seed[2411],seed[1940],seed[1634],seed[117],seed[1565],seed[1025],seed[1172],seed[1720],seed[2274],seed[3660],seed[2299],seed[895],seed[2802],seed[3125],seed[3821],seed[1333],seed[1825],seed[624],seed[3006],seed[3797],seed[1291],seed[2551],seed[492],seed[411],seed[1318],seed[2576],seed[3736],seed[2394],seed[3496],seed[929],seed[903],seed[274],seed[3745],seed[2399],seed[3642],seed[358],seed[2188],seed[1981],seed[3894],seed[120],seed[1788],seed[257],seed[2117],seed[2665],seed[67],seed[3708],seed[1867],seed[3110],seed[3786],seed[2606],seed[601],seed[3123],seed[1506],seed[3492],seed[1273],seed[3883],seed[2888],seed[3068],seed[1950],seed[2482],seed[3377],seed[3101],seed[2890],seed[3257],seed[3678],seed[936],seed[3588],seed[2143],seed[4001],seed[1987],seed[2677],seed[450],seed[2555],seed[2022],seed[3920],seed[683],seed[1659],seed[2466],seed[2945],seed[533],seed[1522],seed[654],seed[2134],seed[3430],seed[2879],seed[2979],seed[3458],seed[1516],seed[865],seed[174],seed[1189],seed[3322],seed[673],seed[1699],seed[632],seed[550],seed[3276],seed[3768],seed[106],seed[820],seed[2430],seed[1780],seed[2041],seed[116],seed[3900],seed[410],seed[2137],seed[2753],seed[2751],seed[9],seed[163],seed[1472],seed[2006],seed[2653],seed[3960],seed[304],seed[288],seed[841],seed[3750],seed[611],seed[551],seed[3511],seed[1602],seed[2846],seed[4060],seed[3399],seed[33],seed[2790],seed[1240],seed[2505],seed[3916],seed[3004],seed[2241],seed[3732],seed[324],seed[1980],seed[811],seed[2773],seed[1875],seed[613],seed[582],seed[3134],seed[1718],seed[3184],seed[1734],seed[3571],seed[1102],seed[3107],seed[536],seed[2726],seed[2974],seed[2807],seed[1731],seed[581],seed[2993],seed[2211],seed[714],seed[3586],seed[2214],seed[334],seed[1035],seed[728],seed[2325],seed[2405],seed[2911],seed[3500],seed[1724],seed[1918],seed[571],seed[1145],seed[3111],seed[1459],seed[3397],seed[405],seed[2320],seed[3555],seed[901],seed[3126],seed[956],seed[1791],seed[2910],seed[2283],seed[2141],seed[3481],seed[3292],seed[3017],seed[4037],seed[1893],seed[2970],seed[112],seed[1892],seed[1941],seed[2581],seed[3159],seed[1443],seed[4061],seed[80],seed[2583],seed[1654],seed[3664],seed[1535],seed[322],seed[3061],seed[3479],seed[604],seed[3537],seed[438],seed[2734],seed[1176],seed[4067],seed[3927],seed[3880],seed[1066],seed[3274],seed[1513],seed[3964],seed[1064],seed[2230],seed[1042],seed[2719],seed[2586],seed[1200],seed[3622],seed[2079],seed[2656],seed[1851],seed[1606],seed[791],seed[4070],seed[840],seed[4003],seed[3728],seed[2179],seed[1316],seed[1835],seed[2874],seed[2617],seed[2454],seed[2263],seed[352],seed[1233],seed[2375],seed[2838],seed[2965],seed[1046],seed[3266],seed[1953],seed[818],seed[2822],seed[63],seed[540],seed[858],seed[346],seed[781],seed[208],seed[1364],seed[425],seed[3790],seed[2703],seed[3130],seed[388],seed[3593],seed[780],seed[3306],seed[3008],seed[2866],seed[1006],seed[2472],seed[2088],seed[923],seed[2172],seed[3164],seed[3902],seed[184],seed[2304],seed[487],seed[3783],seed[483],seed[971],seed[2484],seed[3547],seed[1540],seed[1377],seed[1806],seed[305],seed[31],seed[2836],seed[2308],seed[3684],seed[1763],seed[3007],seed[269],seed[2152],seed[1084],seed[3414],seed[2778],seed[3721],seed[1622],seed[2671],seed[2743],seed[1328],seed[1531],seed[195],seed[3023],seed[453],seed[248],seed[3549],seed[2344],seed[2526],seed[2202],seed[3371],seed[2768],seed[2286],seed[1034],seed[1195],seed[2728],seed[1795],seed[3473],seed[2223],seed[3899],seed[2622],seed[3323],seed[1206],seed[3137],seed[2694],seed[140],seed[938],seed[4044],seed[2765],seed[740],seed[3389],seed[3225],seed[1276],seed[2588],seed[376],seed[480],seed[1792],seed[87],seed[2244],seed[1302],seed[845],seed[1184],seed[463],seed[3962],seed[1394],seed[1842],seed[4084],seed[62],seed[1677],seed[3904],seed[254],seed[386],seed[4074],seed[3709],seed[327],seed[3915],seed[57],seed[761],seed[3602],seed[2389],seed[1614],seed[40],seed[3861],seed[1845],seed[3801],seed[3539],seed[3910],seed[846],seed[860],seed[3752],seed[157],seed[71],seed[264],seed[3887],seed[879],seed[2791],seed[369],seed[3580],seed[3767],seed[1686],seed[23],seed[1451],seed[3772],seed[1434],seed[2412],seed[3143],seed[3019],seed[1804],seed[2135],seed[299],seed[2480],seed[3924],seed[981],seed[690],seed[1905],seed[1674],seed[2207],seed[3975],seed[1714],seed[953],seed[2145],seed[3201],seed[3862],seed[3959],seed[640],seed[298],seed[3109],seed[256],seed[3715],seed[1519],seed[2827],seed[1889],seed[3992],seed[3],seed[24],seed[866],seed[3226],seed[1984],seed[1016],seed[987],seed[3969],seed[3579],seed[3269],seed[1450],seed[105],seed[1109],seed[3616],seed[3097],seed[1815],seed[130],seed[2736],seed[4029],seed[800],seed[441],seed[916],seed[2005],seed[1913],seed[2613],seed[589],seed[1346],seed[996],seed[3273],seed[3365],seed[1124],seed[2563],seed[1169],seed[592],seed[3613],seed[578],seed[1258],seed[1872],seed[1558],seed[2095],seed[2558],seed[3738],seed[394],seed[862],seed[2109],seed[1388],seed[4032],seed[1385],seed[1199],seed[3735],seed[1372],seed[2772],seed[1900],seed[1541],seed[3380],seed[2738],seed[1723],seed[2306],seed[662],seed[1562],seed[2224],seed[3353],seed[2955],seed[3084],seed[1048],seed[2293],seed[716],seed[2718],seed[2545],seed[700],seed[2771],seed[603],seed[3634],seed[995],seed[1611],seed[3546],seed[2146],seed[2165],seed[1221],seed[2075],seed[2932],seed[3319],seed[2410],seed[3394],seed[420],seed[3742],seed[175],seed[3343],seed[736],seed[2462],seed[1164],seed[4049],seed[3597],seed[2056],seed[3015],seed[192],seed[1422],seed[3095],seed[2642],seed[2994],seed[3757],seed[37],seed[2240],seed[3871],seed[1390],seed[2072],seed[4089],seed[4028],seed[3070],seed[1024],seed[4094],seed[1511],seed[3519],seed[2729],seed[1460],seed[2961],seed[3054],seed[1895],seed[2770],seed[3217],seed[287],seed[2784],seed[1678],seed[3596],seed[876],seed[2915],seed[2002],seed[131],seed[1959],seed[460],seed[3557],seed[2739],seed[2854],seed[2083],seed[2478],seed[2654],seed[310],seed[1896],seed[3970],seed[692],seed[1290],seed[827],seed[2914],seed[3648],seed[3706],seed[3698],seed[3753],seed[1742],seed[2196],seed[121],seed[835],seed[775],seed[2535],seed[3466],seed[2851],seed[686],seed[3844],seed[177],seed[2840],seed[4065],seed[1020],seed[3810],seed[1707],seed[1128],seed[2936],seed[2024],seed[1938],seed[3357],seed[1689],seed[2298],seed[1966],seed[2800],seed[717],seed[3946],seed[3552],seed[2052],seed[1823],seed[1452],seed[424],seed[645],seed[1355],seed[788],seed[50],seed[171],seed[3100],seed[2327],seed[2570],seed[445],seed[490],seed[3166],seed[799],seed[1160],seed[147],seed[682],seed[1287],seed[1292],seed[447],seed[1310],seed[366],seed[782],seed[1849],seed[2252],seed[4015],seed[2873],seed[3505],seed[3929],seed[2667],seed[3605],seed[210],seed[56],seed[888],seed[252],seed[529],seed[674],seed[3538],seed[1776],seed[212],seed[1566],seed[3626],seed[2921],seed[2805],seed[241],seed[73],seed[356],seed[349],seed[2939],seed[2826],seed[553],seed[3348],seed[1777],seed[3301],seed[2105],seed[1501],seed[3088],seed[3305],seed[3485],seed[2992],seed[3575],seed[2184],seed[2388],seed[2573],seed[393],seed[1238],seed[3788],seed[3884],seed[3993],seed[3177],seed[3075],seed[3445],seed[3858],seed[1877],seed[594],seed[3621],seed[2003],seed[2107],seed[2036],seed[3467],seed[3132],seed[505],seed[4093],seed[837],seed[558],seed[2102],seed[3477],seed[3944],seed[1770],seed[499],seed[3045],seed[2483],seed[1733],seed[1829],seed[1475],seed[3898],seed[2091],seed[1314],seed[36],seed[2133],seed[3424],seed[2733],seed[68],seed[528],seed[947],seed[3040],seed[3429],seed[1661],seed[2756],seed[3982],seed[30],seed[1473],seed[1616],seed[774],seed[1946],seed[3435],seed[1079],seed[1919],seed[2090],seed[2919],seed[278],seed[1007],seed[684],seed[1901],seed[3565],seed[3014],seed[1643],seed[3791],seed[1843],seed[2029],seed[2725],seed[474],seed[968],seed[99],seed[2000],seed[90],seed[1326],seed[735],seed[2267],seed[1442],seed[2206],seed[2941],seed[2582],seed[1123],seed[2186],seed[778],seed[642],seed[385],seed[2847],seed[1922],seed[235],seed[2457],seed[1440],seed[2301],seed[225],seed[3284],seed[2552],seed[1560],seed[3874],seed[403],seed[17],seed[2048],seed[1487],seed[2812],seed[926],seed[1706],seed[1858],seed[928],seed[2824],seed[198],seed[2780],seed[1075],seed[231],seed[211],seed[3953],seed[3086],seed[2522],seed[3599],seed[951],seed[542],seed[268],seed[3417],seed[833],seed[2931],seed[3703],seed[158],seed[381],seed[4048],seed[21],seed[473],seed[2486],seed[3094],seed[3501],seed[3175],seed[2063],seed[1226],seed[637],seed[1649],seed[4054],seed[2487],seed[2357],seed[2277],seed[1604],seed[2385],seed[3947],seed[1142],seed[2380],seed[100],seed[2110],seed[3631],seed[699],seed[4009],seed[1288],seed[1370],seed[1917],seed[1613],seed[308],seed[3646],seed[185],seed[1332],seed[1635],seed[1219],seed[1975],seed[1995],seed[230],seed[1942],seed[939],seed[3170],seed[3998],seed[671],seed[3794],seed[1873],seed[2549],seed[1568],seed[3345],seed[4010],seed[2816],seed[1642],seed[3295],seed[3923],seed[3199],seed[2130],seed[493],seed[484],seed[3187],seed[2162],seed[564],seed[1876],seed[2720],seed[1651],seed[3326],seed[3216],seed[2721],seed[2348],seed[199],seed[237],seed[11],seed[1340],seed[418],seed[2913],seed[4004],seed[696],seed[896],seed[426],seed[3744],seed[454],seed[917],seed[1054],seed[2010],seed[1799],seed[3531],seed[1929],seed[54],seed[2448],seed[1131],seed[605],seed[580],seed[1805],seed[3643],seed[577],seed[1274],seed[1345],seed[3989],seed[2593],seed[3630],seed[3564],seed[3554],seed[3999],seed[176],seed[78],seed[3667],seed[1703],seed[3925],seed[2132],seed[1347],seed[954],seed[2821],seed[4005],seed[3179],seed[2326],seed[3178],seed[34],seed[1967],seed[3297],seed[164],seed[746],seed[359],seed[3815],seed[2493],seed[1094],seed[1976],seed[3609],seed[1721],seed[357],seed[4038],seed[3160],seed[3193],seed[3892],seed[2111],seed[2958],seed[2875],seed[3259],seed[1391],seed[812],seed[2541],seed[2422],seed[2598],seed[2519],seed[687],seed[3263],seed[576],seed[1914],seed[440],seed[1118],seed[282],seed[317],seed[1790],seed[2343],seed[2722],seed[3651],seed[3085],seed[408],seed[1045],seed[3158],seed[1309],seed[3504],seed[2981],seed[3935],seed[221],seed[732],seed[518],seed[935],seed[3033],seed[3905],seed[3482],seed[2297],seed[1537],seed[2311],seed[1003],seed[1293],seed[3842],seed[1115],seed[3516],seed[2011],seed[1961],seed[597],seed[3229],seed[2391],seed[545],seed[2154],seed[2068],seed[3346],seed[2247],seed[1474],seed[2692],seed[1585],seed[2333],seed[2705],seed[1814],seed[3456],seed[1259],seed[2757],seed[650],seed[88],seed[2216],seed[396],seed[1526],seed[3197],seed[952],seed[4017],seed[1467],seed[2307],seed[2697],seed[20],seed[3816],seed[2521],seed[2354],seed[2349],seed[2264],seed[3053],seed[2950],seed[1486],seed[3120],seed[2167],seed[1068],seed[4045],seed[517],seed[2525],seed[1187],seed[1605],seed[2149],seed[2985],seed[806],seed[1281],seed[2103],seed[2611],seed[3583],seed[2323],seed[3401],seed[364],seed[579],seed[1190],seed[2712],seed[1997],seed[755],seed[1750],seed[69],seed[370],seed[697],seed[3945],seed[3682],seed[569],seed[1878],seed[3455],seed[1081],seed[3983],seed[1228],seed[2225],seed[2023],seed[688],seed[4064],seed[565],seed[3776],seed[253],seed[4025],seed[2131],seed[1303],seed[1725],seed[1523],seed[3612],seed[520],seed[2600],seed[817],seed[3129],seed[2312],seed[678],seed[863],seed[1949],seed[1818],seed[659],seed[368],seed[3432],seed[512],seed[1621],seed[3584],seed[2536],seed[1789],seed[2395],seed[3215],seed[404],seed[3029],seed[2201],seed[1772],seed[306],seed[2474],seed[2151],seed[3627],seed[1671],seed[1225],seed[3113],seed[670],seed[3876],seed[391],seed[667],seed[2446],seed[1398],seed[4091],seed[2066],seed[760],seed[552],seed[2627],seed[2044],seed[2419],seed[3921],seed[1307],seed[3878],seed[2317],seed[267],seed[918],seed[1134],seed[1116],seed[1569],seed[2035],seed[326],seed[1396],seed[3831],seed[1483],seed[3869],seed[3840],seed[1666],seed[871],seed[2749],seed[1193],seed[1402],seed[3384],seed[2129],seed[2537],seed[126],seed[223],seed[2042],seed[3050],seed[10],seed[877],seed[851],seed[295],seed[2510],seed[2475],seed[867],seed[2833],seed[2261],seed[154],seed[4053],seed[949],seed[1751],seed[766],seed[3036],seed[3641],seed[1880],seed[1361],seed[3737],seed[3963],seed[3065],seed[2695],seed[531],seed[2513],seed[1758],seed[2335],seed[2099],seed[1599],seed[2516],seed[2876],seed[3572],seed[2880],seed[1061],seed[1834],seed[749],seed[653],seed[2820],seed[1137],seed[2440],seed[502],seed[3679],seed[1740],seed[2212],seed[1496],seed[1076],seed[839],seed[2946],seed[3051],seed[3800],seed[934],seed[2848],seed[664],seed[1548],seed[1920],seed[514],seed[2696],seed[3202],seed[2465],seed[1538],seed[1080],seed[2124],seed[390],seed[1673],seed[1356],seed[1550],seed[4039],seed[1580],seed[494],seed[2886],seed[1738],seed[1485],seed[1809],seed[789],seed[2358],seed[2810],seed[854],seed[465],seed[1767],seed[2912],seed[2796],seed[2612],seed[1209],seed[1433],seed[1058],seed[1146],seed[2561],seed[2639],seed[1023],seed[629],seed[150],seed[2101],seed[3241],seed[1907],seed[2683],seed[3071],seed[3207],seed[2019],seed[2923],seed[3280],seed[3037],seed[983],seed[1185],seed[3089],seed[899],seed[3524],seed[1037],seed[161],seed[1525],seed[3918],seed[2017],seed[993],seed[2222],seed[111],seed[179],seed[2020],seed[3031],seed[615],seed[1754],seed[2026],seed[1267],seed[2271],seed[219],seed[2907],seed[3696],seed[3867],seed[3663],seed[2530],seed[98],seed[2269],seed[2495],seed[2862],seed[707],seed[2659],seed[3615],seed[181],seed[442],seed[1898],seed[1150],seed[1624],seed[64],seed[1684],seed[2591],seed[1775],seed[3676],seed[3873],seed[1337],seed[340],seed[3282],seed[3073],seed[2776],seed[537],seed[413],seed[2213],seed[1985],seed[3079],seed[2021],seed[2147],seed[1581],seed[1676],seed[906],seed[337],seed[880],seed[94],seed[3337],seed[1234],seed[3958],seed[2903],seed[1968],seed[3623],seed[162],seed[1832],seed[3830],seed[2262],seed[3192],seed[1639],seed[1354],seed[1375],seed[3769],seed[3639],seed[777],seed[3270],seed[2808],seed[2159],seed[1533],seed[1223],seed[259],seed[2996],seed[3152],seed[2782],seed[1557],seed[2741],seed[3145],seed[65],seed[3859],seed[351],seed[3043],seed[205],seed[1021],seed[1295],seed[1904],seed[2787],seed[3055],seed[1435],seed[3581],seed[2603],seed[3324],seed[2938],seed[988],seed[4042],seed[3335],seed[3881],seed[3624],seed[3758],seed[1490],seed[2086],seed[1005],seed[1425],seed[1728],seed[3534],seed[1389],seed[61],seed[2361],seed[3591],seed[3453],seed[2100],seed[2421],seed[3312],seed[372],seed[727],seed[1826],seed[2646],seed[2473],seed[3489],seed[2174],seed[47],seed[1341],seed[1713],seed[4051],seed[665],seed[2070],seed[486],seed[1881],seed[792],seed[965],seed[2713],seed[3955],seed[1050],seed[2497],seed[436],seed[2334],seed[1018],seed[2393],seed[2458],seed[255],seed[3601],seed[3979],seed[2518],seed[753],seed[284],seed[4035],seed[3544],seed[448],seed[821],seed[3025],seed[509],seed[1366],seed[1494],seed[417],seed[3483],seed[3817],seed[427],seed[618],seed[3299],seed[1800],seed[374],seed[1028],seed[320],seed[1479],seed[631],seed[655],seed[1382],seed[3700],seed[280],seed[853],seed[28],seed[1499],seed[1640],seed[893],seed[1685],seed[3978],seed[1521],seed[1194],seed[1837],seed[1426],seed[784],seed[1218],seed[1343],seed[2128],seed[2367],seed[3153],seed[3291],seed[3072],seed[3705],seed[2899],seed[1737],seed[3460],seed[229],seed[2717],seed[3009],seed[2455],seed[2856],seed[1013],seed[2850],seed[2084],seed[2640],seed[2998],seed[2973],seed[977],seed[2256],seed[495],seed[1498],seed[1149],seed[960],seed[770],seed[1031],seed[3361],seed[389],seed[3122],seed[1983],seed[251],seed[3826],seed[2284],seed[2183],seed[1693],seed[4],seed[314],seed[829],seed[1381],seed[1598],seed[3206],seed[1120],seed[3614],seed[2467],seed[1026],seed[1570],seed[414],seed[567],seed[1047],seed[3387],seed[2046],seed[1386],seed[525],seed[2702],seed[2148],seed[3814],seed[1348],seed[2632],seed[354],seed[2935],seed[676],seed[2234],seed[3131],seed[1906],seed[3604],seed[1812],seed[4072],seed[2623],seed[2809],seed[3687],seed[3251],seed[1476],seed[187],seed[3118],seed[3697],seed[718],seed[925],seed[1112],seed[1927],seed[963],seed[3368],seed[2418],seed[1668],seed[1840],seed[3811],seed[2967],seed[3156],seed[1500],seed[2477],seed[4022],seed[3235],seed[872],seed[526],seed[2359],seed[2429],seed[3367],seed[772],seed[530],seed[2924],seed[816],seed[574],seed[3839],seed[1746],seed[1344],seed[1596],seed[3303],seed[661],seed[3330],seed[2877],seed[1441],seed[793],seed[3013],seed[830],seed[2015],seed[2232],seed[290],seed[3162],seed[710],seed[3418],seed[2013],seed[726],seed[294],seed[2673],seed[3710],seed[2715],seed[3124],seed[1785],seed[3294],seed[1179],seed[719],seed[3228],seed[3527],seed[409],seed[3240],seed[1300],seed[2332],seed[997],seed[74],seed[3434],seed[2456],seed[2795],seed[3358],seed[1165],seed[2081],seed[3077],seed[261],seed[962],seed[497],seed[3265],seed[2607],seed[910],seed[1053],seed[2417],seed[123],seed[2698],seed[2315],seed[1629],seed[3403],seed[213],seed[226],seed[713],seed[1368],seed[560],seed[1387],seed[1456],seed[3658],seed[2731],seed[3701],seed[2442],seed[382],seed[1730],seed[2589],seed[3244],seed[992],seed[1682],seed[3933],seed[850],seed[1360],seed[2871],seed[3834],seed[3870],seed[3649],seed[3857],seed[1321],seed[2481],seed[3617],seed[3376],seed[1756],seed[138],seed[3493],seed[2660],seed[2560],seed[3592],seed[2538],seed[1122],seed[3854],seed[4000],seed[1308],seed[1595],seed[3528],seed[1256],seed[331],seed[3115],seed[3606],seed[2173],seed[1862],seed[4095],seed[2089],seed[3942],seed[2533],seed[2777],seed[1732],seed[3359],seed[1552],seed[3069],seed[3940],seed[1033],seed[51],seed[2464],seed[1787],seed[3354],seed[519],seed[3836],seed[606],seed[367],seed[1207],seed[2053],seed[1856],seed[3426],seed[1774],seed[1972],seed[1753],seed[3214],seed[3828],seed[693],seed[908],seed[1888],seed[3675],seed[873],seed[3339],seed[3105],seed[741],seed[489],seed[2381],seed[2595],seed[3363],seed[1],seed[4040],seed[3407],seed[3743],seed[4075],seed[3427],seed[3633],seed[3454],seed[602],seed[643],seed[3587],seed[2450],seed[1235],seed[501],seed[1495],seed[1743],seed[197],seed[2447],seed[1069],seed[3856],seed[3022],seed[2126],seed[3333],seed[1645],seed[2989],seed[4077],seed[3670],seed[946],seed[469],seed[428],seed[737],seed[1726],seed[2832],seed[1493],seed[559],seed[2351],seed[2295],seed[3149],seed[3635],seed[3686],seed[2916],seed[1272],seed[1334],seed[2897],seed[2815],seed[1964],seed[2414],seed[3431],seed[169],seed[1296],seed[1908],seed[2779],seed[3991],seed[2630],seed[2735],seed[3607],seed[3829],seed[842],seed[1930],seed[3808],seed[3535],seed[3749],seed[2038],seed[742],seed[1077],seed[2987],seed[767],seed[3005],seed[986],seed[3136],seed[113],seed[3260],seed[2529],seed[2018],seed[1107],seed[3180],seed[3027],seed[2372],seed[3707],seed[3913],seed[3914],seed[3827],seed[4062],seed[1166],seed[472],seed[1163],seed[3930],seed[2556],seed[344],seed[500],seed[430],seed[360],seed[2905],seed[2409],seed[2532],seed[874],seed[3046],seed[3503],seed[1125],seed[4041],seed[964],seed[2403],seed[620],seed[2187],seed[725],seed[2511],seed[3416],seed[583],seed[58],seed[3347],seed[1482],seed[3433],seed[1974],seed[1484],seed[3780],seed[238],seed[2542],seed[1201],seed[3860],seed[2062],seed[703],seed[1802],seed[244],seed[943],seed[1379],seed[2209],seed[2441],seed[855],seed[1808],seed[466],seed[218],seed[3279],seed[2453],seed[2087],seed[1138],seed[2296],seed[1608],seed[2127],seed[1937],seed[2120],seed[2643],seed[475],seed[3567],seed[1284],seed[1933],seed[2249],seed[1594],seed[1996],seed[193],seed[2275],seed[1220],seed[347],seed[1555],seed[3518],seed[3562],seed[608],seed[2305],seed[824],seed[2723],seed[2892],seed[1576],seed[832],seed[136],seed[375],seed[823],seed[1979],seed[186],seed[1015],seed[3203],seed[109],seed[1641],seed[941],seed[802],seed[155],seed[914],seed[1971],seed[52],seed[3091],seed[456],seed[3719],seed[2689],seed[1764],seed[532],seed[311],seed[554],seed[3994],seed[894],seed[3421],seed[3420],seed[2917],seed[3712],seed[196],seed[3928],seed[3809],seed[2870],seed[3247],seed[3986],seed[160],seed[1264],seed[3603],seed[1243],seed[887],seed[890],seed[128],seed[1263],seed[2788],seed[3973],seed[2428],seed[2944],seed[1119],seed[3486],seed[3001],seed[3314],seed[1289],seed[915],seed[2574],seed[2242],seed[1567],seed[1615],seed[2300],seed[2098],seed[859],seed[82],seed[433],seed[2488],seed[561],seed[1637],seed[3449],seed[214],seed[3837],seed[3666],seed[1374],seed[3764],seed[614],seed[2755],seed[2122],seed[479],seed[808],seed[1657],seed[3931],seed[2266],seed[2631],seed[2259],seed[3150],seed[3480],seed[3852],seed[3689],seed[2553],seed[1087],seed[328],seed[635],seed[2959],seed[1821],seed[2460],seed[745],seed[1988],seed[2814],seed[1405],seed[3230],seed[406],seed[2947],seed[647],seed[1683],seed[3127],seed[292],seed[3315],seed[395],seed[127],seed[2798],seed[1803],seed[1708],seed[12],seed[809],seed[3835],seed[1786],seed[3169],seed[1854],seed[1883],seed[2104],seed[1935],seed[1530],seed[3730],seed[1962],seed[3901],seed[4023],seed[2818],seed[142],seed[3585],seed[3514],seed[429],seed[555],seed[1104],seed[3385],seed[610],seed[1481],seed[1175],seed[3369],seed[1210],seed[2185],seed[2384],seed[4050],seed[89],seed[97],seed[3674],seed[527],seed[1152],seed[3441],seed[1257],seed[2602],seed[1086],seed[2557],seed[1864],seed[1779],seed[151],seed[3632],seed[2675],seed[3509],seed[342],seed[39],seed[658],seed[1097],seed[2064],seed[2074],seed[77],seed[3438],seed[2651],seed[336],seed[3711],seed[1958],seed[146],seed[400],seed[1089],seed[2193],seed[1446],seed[2051],seed[2008],seed[1127],seed[1151],seed[42],seed[3761],seed[4013],seed[2786],seed[3262],seed[1705],seed[4071],seed[731],seed[1099],seed[1191],seed[348],seed[2637],seed[573],seed[2957],seed[2371],seed[2963],seed[3722],seed[2204],seed[139],seed[759],seed[2662],seed[3556],seed[215],seed[2353],seed[1266],seed[1384],seed[1130],seed[4027],seed[621],seed[3714],seed[3655],seed[657],seed[1954],seed[353],seed[1638],seed[2142],seed[3392],seed[3112],seed[3016],seed[2031],seed[3428],seed[3908],seed[4031],seed[4081],seed[1432],seed[3200],seed[1148],seed[2503],seed[1271],seed[2476],seed[3803],seed[3650],seed[590],seed[3465],seed[864],seed[3038],seed[2459],seed[1153],seed[2285],seed[2439],seed[2615],seed[3595],seed[2260],seed[81],seed[1466],seed[630],seed[300],seed[3056],seed[2817],seed[2280],seed[159],seed[3494],seed[2469],seed[3782],seed[1765],seed[3237],seed[2565],seed[932],seed[805],seed[1553],seed[3003],seed[3302],seed[2408],seed[733],seed[1458],seed[3941],seed[3404],seed[3865],seed[2604],seed[764],seed[2281],seed[457],seed[3173],seed[3741],seed[95],seed[3212],seed[2852],seed[3390],seed[2597],seed[3600],seed[3838],seed[1675],seed[2922],seed[3372],seed[2125],seed[1471],seed[321],seed[1010],seed[2071],seed[652],seed[1992],seed[1603],seed[1650],seed[1327],seed[1357],seed[392],seed[1085],seed[2289],seed[1564],seed[398],seed[423],seed[431],seed[1711],seed[1311],seed[1147],seed[4033],seed[1912],seed[1563],seed[144],seed[44],seed[103],seed[2150],seed[3569],seed[3261],seed[3154],seed[3116],seed[2661],seed[521],seed[2057],seed[3488],seed[3798],seed[1952],seed[4080],seed[3440],seed[3577],seed[1245],seed[3720],seed[646],seed[3553],seed[1665],seed[1043],seed[1262],seed[1647],seed[2170],seed[1004],seed[1844],seed[3402],seed[2841],seed[4046],seed[3289],seed[3729],seed[2037],seed[3691],seed[2845],seed[2663],seed[2321],seed[2302],seed[1135],seed[1694],seed[730],seed[3739],seed[3771],seed[2670],seed[838],seed[3598],seed[1229],seed[1820],seed[2716],seed[2272],seed[378],seed[1759],seed[3052],seed[1183],seed[444],seed[3411],seed[4002],seed[467],seed[3227],seed[3298],seed[1978],seed[3396],seed[2507],seed[1982],seed[2085],seed[53],seed[1012],seed[3629],seed[3882],seed[3190],seed[189],seed[974],seed[3476],seed[2766],seed[1778],seed[3672],seed[976],seed[2338],seed[1121],seed[4021],seed[3726],seed[1478],seed[3464],seed[1609],seed[2960],seed[3352],seed[1586],seed[222],seed[2634],seed[1380],seed[2121],seed[539],seed[3032],seed[3618],seed[2254],seed[940],seed[3589],seed[387],seed[2813],seed[283],seed[2363],seed[1994],seed[1508],seed[4069],seed[2392],seed[145],seed[3221],seed[2413],seed[3103],seed[3543],seed[1617],seed[1159],seed[1591],seed[704],seed[1811],seed[2750],seed[3948],seed[2978],seed[644],seed[1692],seed[2547],seed[3926],seed[2709],seed[989],seed[1990],seed[3850],seed[3255],seed[790],seed[2933],seed[3987],seed[758],seed[2370],seed[3340],seed[2452],seed[2045],seed[504],seed[2350],seed[715],seed[1944],seed[249],seed[2954],seed[3189],seed[3802],seed[2584],seed[3774],seed[3787],seed[3657],seed[1891],seed[1002],seed[1957],seed[3172],seed[2164],seed[182],seed[1096],seed[2444],seed[107],seed[137],seed[1866],seed[3886],seed[516],seed[3366],seed[3378],seed[3864],seed[2929],seed[1932],seed[2898],seed[2829],seed[1270],seed[1672],seed[2437],seed[847],seed[1986],seed[1246],seed[984],seed[1539],seed[1108],seed[2055],seed[3762],seed[900],seed[1429],seed[1136],seed[1663],seed[3659],seed[1186],seed[3855],seed[1298],seed[1205],seed[2014],seed[2504],seed[3307],seed[2857],seed[3846],seed[2245],seed[2724],seed[2990],seed[276],seed[762],seed[3082],seed[2679],seed[2449],seed[380],seed[2925],seed[3083],seed[776],seed[1352],seed[102],seed[3512],seed[239],seed[712],seed[1070],seed[3954],seed[1174],seed[470],seed[1378],seed[2889],seed[3747],seed[1860],seed[2764],seed[1633],seed[1871],seed[3563],seed[4066],seed[930],seed[313],seed[2489],seed[1921],seed[3213],seed[702],seed[477],seed[3637],seed[3317],seed[920],seed[1489],seed[148],seed[814],seed[752],seed[2318],seed[570],seed[75],seed[3471],seed[3090],seed[129],seed[1868],seed[3568],seed[2883],seed[2144],seed[118],seed[3288],seed[3640],seed[2839],seed[1943],seed[1143],seed[2969],seed[785],seed[2882],seed[933],seed[399],seed[1524],seed[2198],seed[2984],seed[3796],seed[3042],seed[2253],seed[3231],seed[3695],seed[511],seed[1430],seed[1885],seed[748],seed[2952],seed[2436],seed[1180],seed[156],seed[1559],seed[1410],seed[312],seed[464],seed[1592],seed[2049],seed[1936],seed[1032],seed[705],seed[1027],seed[3048],seed[14],seed[1590],seed[1796],seed[86],seed[3824],seed[1887],seed[3328],seed[416],seed[3047],seed[1545],seed[1114],seed[3239],seed[2975],seed[3452],seed[2789],seed[3521],seed[1749],seed[1991],seed[1359],seed[522],seed[1993],seed[3765],seed[1072],seed[2373],seed[1857],seed[1546],seed[1690],seed[1275],seed[2033],seed[1188],seed[2568],seed[1317],seed[2618],seed[2587],seed[2065],seed[3327],seed[1828],seed[1411],seed[913],seed[1766],seed[3952],seed[1001],seed[663],seed[476],seed[1630],seed[2794],seed[1181],seed[1449],seed[892],seed[978],seed[769],seed[2432],seed[3395],seed[3570],seed[1681],seed[3950],seed[1797],seed[1444],seed[3360],seed[1365],seed[496],seed[3781],seed[3078],seed[3522],seed[641],seed[319],seed[1098],seed[2887],seed[3144],seed[2869],seed[1752],seed[1798],seed[2548],seed[3936],seed[4082],seed[3021],seed[1819],seed[2273],seed[889],seed[1371],seed[544],seed[449],seed[2471],seed[3099],seed[2806],seed[446],seed[3119],seed[1011],seed[1669],seed[3062],seed[596],seed[1505],seed[383],seed[3313],seed[3012],seed[2953],seed[3937],seed[4016],seed[275],seed[3283],seed[3540],seed[1376],seed[3002],seed[1679],seed[2509],seed[166],seed[3000],seed[481],seed[729],seed[2745],seed[2596],seed[2374],seed[2554],seed[919],seed[607],seed[1392],seed[2067],seed[1462],seed[3872],seed[2078],seed[2397],seed[1735],seed[1916],seed[402],seed[471],seed[291],seed[2566],seed[1139],seed[165],seed[91],seed[2175],seed[135],seed[498],seed[1722],seed[3329],seed[1884],seed[1852],seed[2],seed[1008],seed[796],seed[1407],seed[4056],seed[1437],seed[1655],seed[3877],seed[1632],seed[1248],seed[3980],seed[3074],seed[2559],seed[2999],seed[1415],seed[3520],seed[524],seed[2830],seed[3400],seed[3755],seed[1848],seed[85],seed[1232],seed[3063],seed[1626],seed[2027],seed[1126],seed[202],seed[1329],seed[2783],seed[803],seed[508],seed[3995],seed[3219],seed[3717],seed[2398],seed[183],seed[263],seed[2438],seed[2294],seed[1439],seed[3694],seed[4012],seed[3176],seed[309],seed[2161],seed[49],seed[180],seed[1554],seed[458],seed[3891],seed[869],seed[2251],seed[1619],seed[3849],seed[3341],seed[3806],seed[1095],seed[1465],seed[1427],seed[927],seed[4087],seed[2997],seed[27],seed[3997],seed[1251],seed[285],seed[1925],seed[2900],seed[333],seed[3647],seed[343],seed[3264],seed[3656],seed[3704],seed[3690],seed[3139],seed[345],seed[2210],seed[1910],seed[2942],seed[2853],seed[1652],seed[2160],seed[3437],seed[3286],seed[2524],seed[2192],seed[868],seed[1556],seed[191],seed[3813],seed[32],seed[3611],seed[2972],seed[22],seed[4088],seed[622],seed[3669],seed[18],seed[909],seed[2316],seed[739],seed[3141],seed[649],seed[1241],seed[114],seed[1017],seed[2793],seed[891],seed[1306],seed[2415],seed[2215],seed[2620],seed[246],seed[3576],seed[104],seed[2785],seed[3727],seed[1227],seed[373],seed[3102],seed[2759],seed[1762],seed[3406],seed[2097],seed[1768],seed[3066],seed[3943],seed[1561],seed[422],seed[2863],seed[2303],seed[3990],seed[3157],seed[4052],seed[3949],seed[921],seed[3304],seed[2684],seed[4008],seed[1167],seed[2658],seed[844],seed[3868],seed[1544],seed[2178],seed[2649],seed[4011],seed[1036],seed[2629],seed[1280],seed[6],seed[1211],seed[3566],seed[3258],seed[3795],seed[2575],seed[1358],seed[2920],seed[3334],seed[4057],seed[451],seed[3092],seed[1051],seed[1454],seed[1000],seed[273],seed[723],seed[170],seed[3469],seed[1782],seed[3713],seed[2610],seed[3026],seed[1897],seed[2949],seed[1574],seed[3499],seed[751],seed[3638],seed[3243],seed[3041],seed[2693],seed[1696],seed[2203],seed[3785],seed[2106],seed[585],seed[119],seed[70],seed[2616],seed[228],seed[2451],seed[79],seed[355],seed[2747],seed[4079],seed[2331],seed[262],seed[975],seed[3683],seed[3551],seed[3034],seed[2054],seed[1510],seed[1644],seed[3965],seed[1418],seed[1423],seed[1729],seed[3971],seed[3662],seed[3851],seed[2001],seed[3594],seed[260],seed[794],seed[548],seed[3155],seed[1890],seed[3932],seed[1850],seed[1253],seed[1956],seed[216],seed[1784],seed[3423],seed[2878],seed[2569],seed[3491],seed[2797],seed[272],seed[1400],seed[1948],seed[1534],seed[2540],seed[763],seed[2112],seed[1294],seed[681],seed[3773],seed[3128],seed[2191],seed[3236],seed[3804],seed[2231],seed[3723],seed[3560],seed[232],seed[961],seed[2966],seed[3246],seed[3912],seed[2626],seed[3350],seed[2339],seed[1413],seed[3171],seed[1105],seed[2858],seed[303],seed[2140],seed[1573],seed[2523],seed[2276],seed[3974],seed[2199],seed[266],seed[822],seed[595],seed[1299],seed[1547],seed[3412],seed[3439],seed[1453],seed[115],seed[515],seed[861],seed[188],seed[634],seed[2760],seed[2039],seed[970],seed[92],seed[3652],seed[843],seed[297],seed[2156],seed[3985],seed[2943],seed[4076],seed[2257],seed[3351],seed[3383],seed[83],seed[1612],seed[2235],seed[3653],seed[3907],seed[3934],seed[3409],seed[3895],seed[3968],seed[2647],seed[3843],seed[7],seed[1041],seed[3096],seed[1414],seed[2940],seed[1014],seed[134],seed[2636],seed[4036],seed[998],seed[547],seed[4024],seed[1909],seed[96],seed[3956],seed[1970],seed[709],seed[2076],seed[1846],seed[2431],seed[3168],seed[2546],seed[2108],seed[980],seed[810],seed[2073],seed[2435],seed[2976],seed[3463],seed[3897],seed[1646],seed[485],seed[1757],seed[1841],seed[2007],seed[651],seed[1093],seed[1470],seed[1882],seed[2290],seed[125],seed[3725],seed[2287],seed[45],seed[3355],seed[35],seed[1417],seed[2383],seed[3832],seed[3532],seed[1110],seed[3530],seed[2499],seed[2248],seed[1285],seed[2711],seed[2926],seed[990],seed[1648],seed[2605],seed[3415],seed[2706],seed[3718],seed[384],seed[600],seed[3405],seed[3661],seed[2564],seed[307],seed[562],seed[2896],seed[2868],seed[2678],seed[2655],seed[825],seed[1397],seed[3731],seed[924],seed[2506],seed[999],seed[4034],seed[506],seed[3245],seed[1062],seed[1230],seed[1277],seed[2181],seed[2426],seed[1431],seed[3671],seed[1773],seed[4092],seed[1492],seed[4083],seed[459],seed[3805],seed[623],seed[4073],seed[2166],seed[167],seed[379],seed[828],seed[4078],seed[2744],seed[1319],seed[1747],seed[1926],seed[3545],seed[2704],seed[2577],seed[633],seed[362],seed[1588],seed[1101],seed[3468],seed[3507],seed[3558],seed[2842],seed[804],seed[944],seed[3754],seed[3248],seed[3478],seed[982],seed[3349],seed[1171],seed[3451],seed[3370],seed[201],seed[3195],seed[3104],seed[783],seed[826],seed[3939],seed[666],seed[1727],seed[679],seed[3076],seed[1687],seed[2638],seed[1447],seed[549],seed[1260],seed[3853],seed[2685],seed[1618],seed[3142],seed[1320],seed[3256],seed[1448],seed[2329],seed[3194]}),
        .cross_prob(cross_prob),
        .codeword(codeword11),
        .received(received11)
        );
    
    bsc bsc12(
        .clk(clk),
        .reset(reset),
        .seed({seed[1889],seed[3760],seed[1435],seed[3054],seed[2990],seed[3895],seed[1623],seed[3431],seed[1622],seed[3944],seed[1128],seed[2206],seed[3167],seed[3857],seed[2912],seed[1789],seed[215],seed[691],seed[3978],seed[422],seed[957],seed[3940],seed[216],seed[1224],seed[3270],seed[2584],seed[696],seed[3293],seed[1049],seed[322],seed[3074],seed[1216],seed[3135],seed[386],seed[2041],seed[3005],seed[1720],seed[3133],seed[634],seed[1527],seed[2958],seed[2865],seed[2681],seed[966],seed[1436],seed[561],seed[876],seed[2549],seed[37],seed[1201],seed[485],seed[1582],seed[1169],seed[371],seed[301],seed[1648],seed[4002],seed[2062],seed[1108],seed[1865],seed[652],seed[1802],seed[3058],seed[272],seed[2233],seed[3197],seed[2184],seed[1199],seed[580],seed[1034],seed[3141],seed[158],seed[3151],seed[3343],seed[1876],seed[1331],seed[1411],seed[2575],seed[1072],seed[2477],seed[2017],seed[3313],seed[1430],seed[1237],seed[568],seed[1680],seed[2713],seed[3942],seed[1580],seed[665],seed[3998],seed[3236],seed[1280],seed[1801],seed[238],seed[2307],seed[3330],seed[2727],seed[1474],seed[1348],seed[2103],seed[2434],seed[3745],seed[3865],seed[3224],seed[826],seed[3291],seed[3811],seed[708],seed[2904],seed[821],seed[1235],seed[3856],seed[2698],seed[3644],seed[46],seed[2944],seed[1071],seed[4089],seed[2121],seed[3233],seed[2453],seed[3336],seed[3230],seed[2057],seed[1293],seed[3503],seed[2851],seed[1557],seed[401],seed[3273],seed[3264],seed[2197],seed[2693],seed[2910],seed[1499],seed[3189],seed[2678],seed[349],seed[1175],seed[1526],seed[3186],seed[3467],seed[2342],seed[1774],seed[436],seed[3366],seed[3108],seed[2075],seed[2525],seed[2625],seed[551],seed[3458],seed[3098],seed[1185],seed[1406],seed[1251],seed[3],seed[1725],seed[2523],seed[2791],seed[3826],seed[2080],seed[2319],seed[3539],seed[3154],seed[2170],seed[1603],seed[3408],seed[52],seed[1408],seed[2252],seed[889],seed[3164],seed[1518],seed[1891],seed[3551],seed[825],seed[2292],seed[520],seed[2399],seed[2038],seed[1536],seed[563],seed[2669],seed[1573],seed[2978],seed[1200],seed[1521],seed[1964],seed[3365],seed[3424],seed[2995],seed[3119],seed[3850],seed[21],seed[1745],seed[3791],seed[3731],seed[824],seed[2951],seed[3046],seed[2752],seed[4031],seed[521],seed[3742],seed[3908],seed[2943],seed[466],seed[2706],seed[3626],seed[412],seed[359],seed[4077],seed[2209],seed[90],seed[3001],seed[3957],seed[2949],seed[3461],seed[416],seed[2657],seed[1553],seed[290],seed[4039],seed[3795],seed[903],seed[441],seed[1697],seed[885],seed[3331],seed[3451],seed[2831],seed[3816],seed[1424],seed[455],seed[1578],seed[3846],seed[2249],seed[3335],seed[3262],seed[1286],seed[2253],seed[264],seed[2579],seed[2915],seed[3225],seed[3538],seed[2553],seed[1957],seed[3871],seed[60],seed[2665],seed[2235],seed[1857],seed[913],seed[1461],seed[3936],seed[2690],seed[3735],seed[3955],seed[1555],seed[3891],seed[2378],seed[103],seed[1595],seed[3641],seed[294],seed[526],seed[556],seed[2371],seed[2458],seed[3147],seed[2212],seed[245],seed[3199],seed[3642],seed[738],seed[1862],seed[904],seed[527],seed[1630],seed[1088],seed[1830],seed[2231],seed[312],seed[130],seed[395],seed[3607],seed[1223],seed[2430],seed[2815],seed[1144],seed[397],seed[3802],seed[1405],seed[1104],seed[1043],seed[3102],seed[2446],seed[2980],seed[1266],seed[3550],seed[3452],seed[2590],seed[848],seed[1998],seed[2333],seed[1395],seed[763],seed[1033],seed[1698],seed[2177],seed[2269],seed[410],seed[405],seed[2408],seed[3914],seed[2077],seed[3290],seed[2247],seed[2683],seed[4006],seed[263],seed[253],seed[1619],seed[3789],seed[658],seed[92],seed[1315],seed[757],seed[2884],seed[1272],seed[3268],seed[2410],seed[4082],seed[1150],seed[2945],seed[3276],seed[3041],seed[3966],seed[3591],seed[1139],seed[678],seed[991],seed[6],seed[2878],seed[1490],seed[4005],seed[995],seed[4020],seed[3967],seed[3980],seed[2830],seed[1911],seed[469],seed[2517],seed[1361],seed[1123],seed[1805],seed[2747],seed[2519],seed[3706],seed[667],seed[3127],seed[3298],seed[969],seed[2507],seed[370],seed[3606],seed[180],seed[609],seed[2159],seed[3462],seed[1611],seed[2028],seed[1415],seed[1892],seed[554],seed[1429],seed[666],seed[203],seed[3311],seed[4072],seed[91],seed[3316],seed[1218],seed[2597],seed[3919],seed[1585],seed[772],seed[1277],seed[3240],seed[3993],seed[1012],seed[2628],seed[2297],seed[127],seed[449],seed[3410],seed[472],seed[3786],seed[73],seed[417],seed[2711],seed[2930],seed[163],seed[1899],seed[3718],seed[1559],seed[2210],seed[3694],seed[1058],seed[2667],seed[2610],seed[2435],seed[3488],seed[484],seed[3161],seed[523],seed[2604],seed[3571],seed[3960],seed[2006],seed[854],seed[880],seed[1810],seed[1133],seed[3977],seed[2725],seed[599],seed[3125],seed[733],seed[140],seed[2736],seed[2056],seed[3035],seed[3471],seed[3509],seed[3725],seed[861],seed[289],seed[67],seed[3738],seed[3754],seed[3665],seed[1079],seed[1303],seed[2534],seed[898],seed[1860],seed[1078],seed[795],seed[1824],seed[2709],seed[4028],seed[126],seed[1843],seed[3817],seed[593],seed[4015],seed[2989],seed[850],seed[1628],seed[1528],seed[994],seed[1186],seed[2443],seed[2364],seed[2244],seed[4093],seed[1649],seed[2360],seed[2417],seed[1180],seed[3423],seed[2198],seed[2139],seed[11],seed[2708],seed[4085],seed[128],seed[2528],seed[1492],seed[3118],seed[3672],seed[3689],seed[549],seed[1929],seed[25],seed[1846],seed[2465],seed[1909],seed[2536],seed[618],seed[2354],seed[1346],seed[1096],seed[1325],seed[3324],seed[1294],seed[934],seed[204],seed[746],seed[2243],seed[1692],seed[2302],seed[1829],seed[1716],seed[74],seed[547],seed[1941],seed[3958],seed[145],seed[3381],seed[2228],seed[2048],seed[1335],seed[3649],seed[2167],seed[1242],seed[3755],seed[2343],seed[3003],seed[2758],seed[3299],seed[1020],seed[3409],seed[646],seed[1153],seed[2415],seed[1520],seed[2000],seed[1141],seed[3403],seed[1493],seed[85],seed[2969],seed[751],seed[985],seed[482],seed[305],seed[2270],seed[246],seed[1517],seed[2495],seed[684],seed[3188],seed[905],seed[2612],seed[356],seed[232],seed[2763],seed[468],seed[1779],seed[3620],seed[1589],seed[278],seed[2572],seed[1212],seed[4063],seed[3357],seed[835],seed[3628],seed[423],seed[3375],seed[3066],seed[3938],seed[4084],seed[1664],seed[2786],seed[2992],seed[3079],seed[3518],seed[3126],seed[1672],seed[3630],seed[2921],seed[1715],seed[641],seed[2405],seed[149],seed[1906],seed[4035],seed[3068],seed[2149],seed[595],seed[344],seed[1606],seed[292],seed[1481],seed[632],seed[3282],seed[1788],seed[3608],seed[2308],seed[793],seed[2923],seed[3781],seed[3541],seed[884],seed[3281],seed[2986],seed[681],seed[178],seed[385],seed[1885],seed[1130],seed[831],seed[2190],seed[40],seed[376],seed[133],seed[2412],seed[3807],seed[1285],seed[791],seed[2613],seed[1888],seed[1073],seed[2996],seed[944],seed[2794],seed[3542],seed[1412],seed[1060],seed[1665],seed[3612],seed[2275],seed[3679],seed[2259],seed[1143],seed[2451],seed[1349],seed[1304],seed[3768],seed[3269],seed[2288],seed[137],seed[1117],seed[1152],seed[516],seed[10],seed[2508],seed[3783],seed[2471],seed[328],seed[662],seed[2551],seed[2934],seed[2714],seed[1148],seed[3130],seed[1134],seed[3416],seed[3002],seed[477],seed[1399],seed[1605],seed[352],seed[3599],seed[788],seed[1763],seed[2619],seed[1712],seed[853],seed[1897],seed[3711],seed[870],seed[3156],seed[3563],seed[1506],seed[2592],seed[94],seed[2658],seed[3229],seed[2036],seed[2805],seed[3976],seed[142],seed[2386],seed[2457],seed[3194],seed[1807],seed[2656],seed[1693],seed[1917],seed[64],seed[2204],seed[1933],seed[743],seed[2039],seed[1197],seed[1268],seed[2699],seed[3825],seed[3379],seed[1247],seed[1145],seed[1271],seed[3413],seed[175],seed[220],seed[1083],seed[2445],seed[300],seed[132],seed[4062],seed[2882],seed[1187],seed[2467],seed[752],seed[1566],seed[940],seed[2183],seed[1390],seed[3097],seed[768],seed[562],seed[1529],seed[434],seed[2274],seed[1753],seed[62],seed[3279],seed[3842],seed[3243],seed[4040],seed[2131],seed[3866],seed[148],seed[3280],seed[1136],seed[2479],seed[956],seed[1717],seed[2670],seed[1916],seed[3176],seed[1702],seed[1507],seed[3064],seed[2854],seed[2751],seed[3110],seed[34],seed[697],seed[2723],seed[13],seed[2807],seed[3090],seed[465],seed[989],seed[3992],seed[1831],seed[3572],seed[1161],seed[1063],seed[4017],seed[1240],seed[3227],seed[2128],seed[1749],seed[3247],seed[1950],seed[2558],seed[888],seed[3000],seed[1439],seed[2700],seed[14],seed[2361],seed[3892],seed[1385],seed[3534],seed[2540],seed[3592],seed[2810],seed[2648],seed[1784],seed[2340],seed[2710],seed[2685],seed[740],seed[700],seed[3007],seed[571],seed[1082],seed[3870],seed[3323],seed[1051],seed[1598],seed[3426],seed[1848],seed[2491],seed[491],seed[2188],seed[637],seed[2724],seed[1524],seed[1669],seed[2223],seed[2050],seed[922],seed[4049],seed[2054],seed[297],seed[3882],seed[1711],seed[1444],seed[3078],seed[1227],seed[1983],seed[1232],seed[1539],seed[2439],seed[1639],seed[1990],seed[1821],seed[1914],seed[2022],seed[3739],seed[1509],seed[2127],seed[3748],seed[1599],seed[3277],seed[3080],seed[2178],seed[155],seed[2639],seed[1334],seed[1228],seed[2239],seed[2950],seed[3433],seed[3506],seed[1770],seed[2413],seed[3660],seed[654],seed[2688],seed[3931],seed[1955],seed[924],seed[820],seed[660],seed[3762],seed[1151],seed[3838],seed[2746],seed[3449],seed[2858],seed[2749],seed[2225],seed[4007],seed[1650],seed[467],seed[265],seed[3310],seed[2643],seed[965],seed[2011],seed[348],seed[3872],seed[745],seed[440],seed[3180],seed[2119],seed[3740],seed[3564],seed[3831],seed[343],seed[1569],seed[3082],seed[2144],seed[1695],seed[2448],seed[3019],seed[3470],seed[3637],seed[1744],seed[1627],seed[3474],seed[1996],seed[2913],seed[1262],seed[2888],seed[4019],seed[2599],seed[3445],seed[2407],seed[4034],seed[2087],seed[1236],seed[439],seed[2899],seed[3190],seed[1155],seed[2767],seed[2580],seed[2004],seed[2273],seed[3201],seed[3686],seed[2973],seed[3393],seed[570],seed[2015],seed[286],seed[584],seed[1596],seed[86],seed[2661],seed[1505],seed[3521],seed[711],seed[2102],seed[926],seed[3105],seed[972],seed[3034],seed[2256],seed[2304],seed[2433],seed[642],seed[3692],seed[45],seed[2023],seed[2692],seed[1985],seed[3766],seed[1905],seed[4080],seed[3528],seed[239],seed[2979],seed[4087],seed[1718],seed[1039],seed[3851],seed[2179],seed[494],seed[1401],seed[2780],seed[3926],seed[1122],seed[3884],seed[28],seed[897],seed[3578],seed[2920],seed[2005],seed[2328],seed[1340],seed[3049],seed[3537],seed[1626],seed[1095],seed[2608],seed[1781],seed[3193],seed[2109],seed[3719],seed[2030],seed[1523],seed[4073],seed[374],seed[535],seed[2373],seed[2897],seed[3833],seed[1026],seed[921],seed[2353],seed[1875],seed[3439],seed[3670],seed[3255],seed[2679],seed[935],seed[2018],seed[2376],seed[907],seed[3380],seed[2146],seed[1867],seed[2151],seed[1577],seed[3505],seed[2538],seed[3008],seed[110],seed[1488],seed[3805],seed[1545],seed[2444],seed[1561],seed[2120],seed[3210],seed[805],seed[3587],seed[3604],seed[3140],seed[2002],seed[727],seed[776],seed[2012],seed[2855],seed[1618],seed[3484],seed[1011],seed[3138],seed[1061],seed[1683],seed[2403],seed[3177],seed[1609],seed[2676],seed[1567],seed[1485],seed[497],seed[1041],seed[3069],seed[219],seed[1306],seed[3533],seed[1471],seed[3249],seed[2324],seed[458],seed[2492],seed[2694],seed[2089],seed[2909],seed[674],seed[167],seed[3038],seed[685],seed[3317],seed[933],seed[3026],seed[3989],seed[3737],seed[3651],seed[1883],seed[1930],seed[2890],seed[2073],seed[2626],seed[1312],seed[2422],seed[4004],seed[742],seed[3139],seed[760],seed[1548],seed[1787],seed[4044],seed[1313],seed[3655],seed[1961],seed[2152],seed[582],seed[3212],seed[3894],seed[3522],seed[895],seed[2115],seed[1057],seed[2021],seed[699],seed[1383],seed[1069],seed[2938],seed[1615],seed[3513],seed[2808],seed[669],seed[3111],seed[2594],seed[1901],seed[2],seed[1065],seed[2175],seed[3800],seed[3921],seed[1834],seed[3812],seed[1419],seed[2141],seed[592],seed[65],seed[2889],seed[2772],seed[2192],seed[3773],seed[3460],seed[1179],seed[2091],seed[1847],seed[2860],seed[3981],seed[2086],seed[1105],seed[29],seed[1602],seed[1106],seed[1691],seed[3367],seed[838],seed[1912],seed[2903],seed[27],seed[3621],seed[2827],seed[1341],seed[3114],seed[197],seed[3036],seed[460],seed[53],seed[533],seed[3923],seed[2722],seed[1017],seed[651],seed[2045],seed[3574],seed[3619],seed[3830],seed[3368],seed[1854],seed[2589],seed[3887],seed[3517],seed[522],seed[3597],seed[3933],seed[2695],seed[2562],seed[544],seed[256],seed[2305],seed[873],seed[1965],seed[1070],seed[1050],seed[1962],seed[2291],seed[2524],seed[2646],seed[2790],seed[2416],seed[190],seed[1005],seed[3319],seed[87],seed[3788],seed[1167],seed[815],seed[1554],seed[3158],seed[1677],seed[2237],seed[3615],seed[2485],seed[4067],seed[1337],seed[1953],seed[251],seed[1489],seed[2287],seed[2922],seed[3687],seed[529],seed[2759],seed[3875],seed[2497],seed[1927],seed[2985],seed[2647],seed[3456],seed[910],seed[2891],seed[3198],seed[892],seed[2964],seed[877],seed[3347],seed[2129],seed[2147],seed[2272],seed[2875],seed[3581],seed[1336],seed[611],seed[2455],seed[315],seed[2828],seed[1426],seed[2629],seed[2166],seed[3526],seed[2998],seed[1465],seed[61],seed[2777],seed[2283],seed[2560],seed[4074],seed[336],seed[1794],seed[1920],seed[2935],seed[3106],seed[1999],seed[3569],seed[2164],seed[3954],seed[1098],seed[3245],seed[1413],seed[2853],seed[369],seed[605],seed[2258],seed[3968],seed[1607],seed[1015],seed[1844],seed[1475],seed[1160],seed[3639],seed[2122],seed[2573],seed[41],seed[3478],seed[3720],seed[3053],seed[3905],seed[3318],seed[1305],seed[602],seed[2230],seed[3710],seed[655],seed[3787],seed[3705],seed[75],seed[616],seed[1328],seed[1783],seed[3836],seed[1101],seed[1456],seed[3314],seed[2196],seed[3004],seed[581],seed[3132],seed[3983],seed[3344],seed[2529],seed[2049],seed[229],seed[196],seed[3784],seed[420],seed[714],seed[836],seed[589],seed[1460],seed[2401],seed[3271],seed[66],seed[392],seed[3417],seed[799],seed[3384],seed[2662],seed[3415],seed[2263],seed[1402],seed[607],seed[247],seed[875],seed[2363],seed[1410],seed[2173],seed[623],seed[1149],seed[560],seed[47],seed[1102],seed[3822],seed[213],seed[1124],seed[2511],seed[3829],seed[3283],seed[3429],seed[1332],seed[649],seed[1931],seed[3045],seed[2927],seed[483],seed[2718],seed[868],seed[3308],seed[3399],seed[3839],seed[1678],seed[2214],seed[1719],seed[1841],seed[2883],seed[2817],seed[3202],seed[2555],seed[235],seed[2500],seed[172],seed[1881],seed[3238],seed[2279],seed[2541],seed[2505],seed[381],seed[1737],seed[3371],seed[3163],seed[1740],seed[3124],seed[2462],seed[950],seed[4051],seed[1296],seed[1183],seed[2241],seed[1252],seed[578],seed[2499],seed[4056],seed[1154],seed[273],seed[3912],seed[997],seed[150],seed[1202],seed[2917],seed[3434],seed[1255],seed[3083],seed[2084],seed[1441],seed[1035],seed[16],seed[983],seed[2418],seed[1519],seed[753],seed[1706],seed[1747],seed[368],seed[3761],seed[628],seed[2717],seed[871],seed[3500],seed[2929],seed[1945],seed[3267],seed[1701],seed[3376],seed[778],seed[722],seed[729],seed[2602],seed[4030],seed[3752],seed[3614],seed[594],seed[2886],seed[3671],seed[2901],seed[2208],seed[3169],seed[2754],seed[3350],seed[1068],seed[3730],seed[1882],seed[327],seed[2171],seed[785],seed[364],seed[20],seed[354],seed[4066],seed[1771],seed[2850],seed[3244],seed[3510],seed[144],seed[1376],seed[459],seed[3749],seed[451],seed[1416],seed[1014],seed[1915],seed[3094],seed[900],seed[786],seed[998],seed[100],seed[917],seed[1730],seed[3662],seed[1244],seed[2741],seed[2587],seed[489],seed[2372],seed[2298],seed[971],seed[4033],seed[2906],seed[928],seed[32],seed[2680],seed[1635],seed[3285],seed[230],seed[3585],seed[967],seed[2892],seed[902],seed[683],seed[307],seed[3855],seed[2156],seed[2470],seed[1168],seed[2282],seed[3454],seed[3172],seed[1006],seed[2172],seed[2516],seed[3516],seed[3485],seed[329],seed[1100],seed[908],seed[3329],seed[932],seed[2161],seed[139],seed[225],seed[4003],seed[1194],seed[3514],seed[1283],seed[2421],seed[3191],seed[2863],seed[1044],seed[1856],seed[1319],seed[3187],seed[4053],seed[1726],seed[1560],seed[310],seed[3647],seed[3373],seed[2094],seed[878],seed[1658],seed[1647],seed[3849],seed[182],seed[1594],seed[2406],seed[1620],seed[3322],seed[591],seed[1780],seed[3301],seed[3061],seed[704],seed[1025],seed[2357],seed[3498],seed[4050],seed[165],seed[3144],seed[1919],seed[4069],seed[268],seed[2707],seed[3043],seed[1980],seed[2644],seed[503],seed[1177],seed[3906],seed[1657],seed[3013],seed[3907],seed[3383],seed[2814],seed[226],seed[2955],seed[2180],seed[866],seed[2150],seed[942],seed[107],seed[1275],seed[3683],seed[2490],seed[2849],seed[2874],seed[1380],seed[915],seed[379],seed[1323],seed[2653],seed[1835],seed[2398],seed[961],seed[2603],seed[2240],seed[3530],seed[2303],seed[2033],seed[2003],seed[2313],seed[726],seed[2436],seed[3899],seed[2804],seed[3600],seed[576],seed[3214],seed[1450],seed[2203],seed[1687],seed[1090],seed[314],seed[2227],seed[2383],seed[83],seed[1353],seed[3820],seed[883],seed[2392],seed[1250],seed[3185],seed[2125],seed[1084],seed[2459],seed[3305],seed[3814],seed[1066],seed[3951],seed[1676],seed[672],seed[181],seed[698],seed[695],seed[1320],seed[3407],seed[3877],seed[3724],seed[2545],seed[1491],seed[3927],seed[3668],seed[1024],seed[1116],seed[3646],seed[2556],seed[511],seed[1081],seed[193],seed[138],seed[1111],seed[1616],seed[688],seed[1816],seed[3042],seed[2079],seed[1270],seed[2994],seed[2182],seed[1799],seed[1156],seed[2836],seed[3442],seed[2309],seed[759],seed[2335],seed[1951],seed[1479],seed[3237],seed[1302],seed[2800],seed[1734],seed[1356],seed[1671],seed[4047],seed[2290],seed[3695],seed[2673],seed[345],seed[63],seed[316],seed[1790],seed[1219],seed[1866],seed[3022],seed[920],seed[3027],seed[2503],seed[2099],seed[2654],seed[357],seed[1056],seed[3494],seed[762],seed[2637],seed[3726],seed[719],seed[214],seed[2677],seed[758],seed[2702],seed[3501],seed[3047],seed[1689],seed[3904],seed[1099],seed[2965],seed[1796],seed[1495],seed[2068],seed[3203],seed[4026],seed[1913],seed[1478],seed[2327],seed[3939],seed[3536],seed[1572],seed[1637],seed[1604],seed[811],seed[1556],seed[1873],seed[2696],seed[1688],seed[3263],seed[2916],seed[2861],seed[3840],seed[2911],seed[2475],seed[2820],seed[3174],seed[2729],seed[3780],seed[2472],seed[2261],seed[2163],seed[679],seed[1085],seed[1574],seed[2788],seed[1670],seed[1038],seed[1046],seed[675],seed[3885],seed[174],seed[510],seed[3828],seed[525],seed[3075],seed[2034],seed[781],seed[1022],seed[1516],seed[2530],seed[3702],seed[1995],seed[112],seed[1103],seed[2266],seed[114],seed[1992],seed[555],seed[2900],seed[2796],seed[1721],seed[960],seed[2756],seed[1273],seed[1817],seed[54],seed[3696],seed[3965],seed[2601],seed[566],seed[1513],seed[1284],seed[718],seed[1254],seed[702],seed[1295],seed[1203],seed[2104],seed[2348],seed[4012],seed[2130],seed[1003],seed[1125],seed[955],seed[3941],seed[2778],seed[3120],seed[3428],seed[1758],seed[2847],seed[689],seed[1469],seed[3232],seed[1984],seed[2533],seed[492],seed[1394],seed[1459],seed[2154],seed[2118],seed[2504],seed[3909],seed[659],seed[865],seed[744],seed[2844],seed[1354],seed[3974],seed[1409],seed[1925],seed[173],seed[993],seed[3476],seed[3611],seed[3018],seed[3845],seed[2420],seed[862],seed[919],seed[81],seed[3512],seed[2277],seed[1274],seed[1500],seed[1008],seed[2058],seed[860],seed[2856],seed[2873],seed[3582],seed[478],seed[1837],seed[129],seed[2264],seed[3101],seed[3360],seed[2789],seed[3395],seed[2926],seed[2521],seed[3136],seed[1142],seed[1887],seed[2512],seed[341],seed[2947],seed[3535],seed[1427],seed[1923],seed[2318],seed[1993],seed[1301],seed[2582],seed[3205],seed[1486],seed[2840],seed[3547],seed[2138],seed[2338],seed[3063],seed[51],seed[481],seed[1870],seed[2832],seed[3231],seed[3432],seed[1448],seed[1338],seed[687],seed[3767],seed[2060],seed[2400],seed[3020],seed[1926],seed[339],seed[4083],seed[3014],seed[3540],seed[822],seed[2771],seed[1575],seed[1979],seed[946],seed[2928],seed[1540],seed[3774],seed[1772],seed[2755],seed[3195],seed[2715],seed[400],seed[1404],seed[1714],seed[1989],seed[622],seed[2114],seed[2531],seed[2052],seed[453],seed[1037],seed[1166],seed[4029],seed[2143],seed[1674],seed[1681],seed[3048],seed[4070],seed[3583],seed[3307],seed[136],seed[1551],seed[1633],seed[378],seed[2966],seed[1751],seed[3779],seed[2522],seed[775],seed[1853],seed[627],seed[1795],seed[1653],seed[2332],seed[2195],seed[810],seed[615],seed[3995],seed[1047],seed[3584],seed[3295],seed[2255],seed[677],seed[3853],seed[3697],seed[4032],seed[38],seed[2615],seed[604],seed[1700],seed[2569],seed[3799],seed[2846],seed[2137],seed[1601],seed[1019],seed[620],seed[212],seed[210],seed[430],seed[121],seed[2914],seed[2098],seed[2552],seed[930],seed[280],seed[1898],seed[4048],seed[3459],seed[2450],seed[970],seed[108],seed[2869],seed[703],seed[2887],seed[1453],seed[2671],seed[3673],seed[3677],seed[3502],seed[2720],seed[3848],seed[518],seed[2359],seed[3753],seed[1221],seed[2801],seed[1207],seed[650],seed[1198],seed[818],seed[890],seed[118],seed[1921],seed[1769],seed[3148],seed[1852],seed[452],seed[1355],seed[2879],seed[3491],seed[1428],seed[2982],seed[3477],seed[1684],seed[160],seed[1591],seed[3093],seed[3463],seed[2924],seed[2339],seed[725],seed[1174],seed[2201],seed[2019],seed[1109],seed[852],seed[3032],seed[1859],seed[1818],seed[1703],seed[1510],seed[4013],seed[1278],seed[2806],seed[3159],seed[3055],seed[1241],seed[574],seed[285],seed[2781],seed[857],seed[279],seed[2219],seed[2257],seed[3804],seed[546],seed[539],seed[3192],seed[2750],seed[625],seed[3143],seed[1327],seed[415],seed[1009],seed[1625],seed[806],seed[1466],seed[1825],seed[4022],seed[3059],seed[567],seed[737],seed[626],seed[1590],seed[2107],seed[1127],seed[1632],seed[1982],seed[2775],seed[2007],seed[2390],seed[978],seed[323],seed[3092],seed[2894],seed[1994],seed[664],seed[3910],seed[3328],seed[3810],seed[2797],seed[84],seed[1021],seed[3402],seed[1359],seed[3801],seed[1248],seed[1414],seed[4046],seed[572],seed[864],seed[3364],seed[927],seed[2967],seed[3123],seed[2730],seed[3396],seed[396],seed[1075],seed[2194],seed[3566],seed[3699],seed[2682],seed[1814],seed[1205],seed[1791],seed[528],seed[2218],seed[3529],seed[260],seed[2632],seed[3028],seed[2948],seed[2145],seed[2812],seed[170],seed[3782],seed[1059],seed[1324],seed[3721],seed[2111],seed[1798],seed[2616],seed[1129],seed[701],seed[2396],seed[366],seed[1292],seed[977],seed[2083],seed[2042],seed[3287],seed[3504],seed[2867],seed[97],seed[2330],seed[2954],seed[1132],seed[3024],seed[3346],seed[3015],seed[2997],seed[1537],seed[1114],seed[2585],seed[918],seed[2380],seed[3631],seed[1903],seed[2454],seed[2460],seed[1864],seed[2704],seed[3656],seed[1833],seed[519],seed[2064],seed[517],seed[2893],seed[954],seed[1172],seed[3216],seed[1958],seed[332],seed[3349],seed[1112],seed[3924],seed[1115],seed[2957],seed[9],seed[2548],seed[1352],seed[346],seed[588],seed[3854],seed[244],seed[2488],seed[2550],seed[2798],seed[2618],seed[388],seed[179],seed[715],seed[373],seed[851],seed[3765],seed[779],seed[3095],seed[143],seed[2423],seed[721],seed[3837],seed[1329],seed[3552],seed[3261],seed[1952],seed[807],seed[1000],seed[3969],seed[1501],seed[2737],seed[1029],seed[77],seed[2481],seed[2323],seed[657],seed[1027],seed[2535],seed[1742],seed[33],seed[1815],seed[313],seed[1372],seed[2649],seed[4052],seed[1403],seed[887],seed[2331],seed[1288],seed[847],seed[2976],seed[406],seed[735],seed[1291],seed[456],seed[1690],seed[3217],seed[3573],seed[630],seed[269],seed[512],seed[2566],seed[2486],seed[1662],seed[2933],seed[3827],seed[3052],seed[2306],seed[4065],seed[2848],seed[4095],seed[2953],seed[3580],seed[1785],seed[30],seed[1624],seed[1544],seed[2666],seed[281],seed[2334],seed[3863],seed[199],seed[3181],seed[717],seed[1362],seed[1813],seed[3729],seed[841],seed[3627],seed[1682],seed[1384],seed[1822],seed[1535],seed[1257],seed[2296],seed[2735],seed[1258],seed[3691],seed[487],seed[790],seed[2972],seed[1502],seed[2547],seed[1373],seed[4009],seed[3722],seed[2742],seed[3325],seed[2819],seed[3684],seed[258],seed[564],seed[769],seed[43],seed[1126],seed[1016],seed[147],seed[1872],seed[19],seed[2782],seed[2356],seed[1565],seed[2464],seed[2761],seed[1253],seed[3128],seed[1608],seed[3618],seed[710],seed[3170],seed[2326],seed[2397],seed[3253],seed[1515],seed[3970],seed[2097],seed[3129],seed[794],seed[2440],seed[1457],seed[3497],seed[2384],seed[3440],seed[3254],seed[2574],seed[1863],seed[3868],seed[1991],seed[1970],seed[557],seed[1454],seed[2375],seed[540],seed[1612],seed[2478],seed[3411],seed[2543],seed[2442],seed[2870],seed[1091],seed[454],seed[3387],seed[3222],seed[3011],seed[1651],seed[1543],seed[3259],seed[168],seed[2857],seed[284],seed[2532],seed[1773],seed[3398],seed[2250],seed[186],seed[3418],seed[3985],seed[1724],seed[1417],seed[2135],seed[819],seed[464],seed[3678],seed[261],seed[399],seed[1775],seed[748],seed[1196],seed[2293],seed[1163],seed[3178],seed[241],seed[1443],seed[1811],seed[351],seed[404],seed[2544],seed[1778],seed[1571],seed[3950],seed[1287],seed[3242],seed[486],seed[96],seed[1260],seed[3659],seed[796],seed[2672],seed[2238],seed[3664],seed[1842],seed[4038],seed[1269],seed[3303],seed[2321],seed[78],seed[3115],seed[2085],seed[3155],seed[893],seed[48],seed[3466],seed[4042],seed[1425],seed[473],seed[2320],seed[1954],seed[712],seed[1389],seed[293],seed[3397],seed[1229],seed[3532],seed[2770],seed[899],seed[2093],seed[324],seed[2126],seed[541],seed[3545],seed[350],seed[986],seed[1878],seed[4008],seed[937],seed[2902],seed[923],seed[1377],seed[1256],seed[739],seed[3511],seed[1549],seed[783],seed[2301],seed[2743],seed[3771],seed[298],seed[2369],seed[1358],seed[3523],seed[3033],seed[499],seed[228],seed[3081],seed[1318],seed[1968],seed[2636],seed[3548],seed[1819],seed[1673],seed[1300],seed[680],seed[3629],seed[2381],seed[645],seed[3208],seed[2593],seed[3878],seed[1189],seed[1476],seed[1849],seed[1765],seed[1708],seed[131],seed[2035],seed[4037],seed[335],seed[3727],seed[3312],seed[610],seed[3815],seed[3386],seed[2082],seed[2826],seed[3076],seed[3337],seed[55],seed[2962],seed[803],seed[1587],seed[1210],seed[218],seed[2113],seed[3930],seed[2687],seed[1363],seed[2631],seed[2689],seed[1894],seed[1886],seed[1146],seed[377],seed[3309],seed[2181],seed[2868],seed[3601],seed[479],seed[509],seed[1048],seed[736],seed[3712],seed[1729],seed[3893],seed[988],seed[2939],seed[4018],seed[916],seed[2176],seed[3131],seed[2627],seed[2960],seed[1370],seed[488],seed[2617],seed[545],seed[2838],seed[1826],seed[3029],seed[614],seed[1614],seed[2026],seed[1741],seed[2200],seed[187],seed[1550],seed[827],seed[367],seed[3107],seed[1757],seed[1093],seed[3949],seed[200],seed[3874],seed[3218],seed[2385],seed[363],seed[421],seed[382],seed[3746],seed[2956],seed[2809],seed[3700],seed[387],seed[3602],seed[3353],seed[2222],seed[2701],seed[947],seed[3362],seed[1646],seed[2557],seed[3252],seed[2047],seed[2009],seed[3759],seed[217],seed[814],seed[2784],seed[2799],seed[3358],seed[2031],seed[1710],seed[2931],seed[437],seed[2216],seed[1067],seed[2919],seed[943],seed[797],seed[1137],seed[2576],seed[2732],seed[70],seed[3775],seed[360],seed[798],seed[912],seed[4010],seed[3717],seed[756],seed[3257],seed[3040],seed[3378],seed[471],seed[2733],seed[1343],seed[3603],seed[240],seed[3184],seed[2136],seed[4058],seed[2765],seed[3867],seed[843],seed[728],seed[2351],seed[1694],seed[3888],seed[361],seed[1445],seed[3421],seed[3847],seed[3294],seed[1282],seed[1823],seed[1713],seed[3085],seed[3616],seed[2651],seed[2981],seed[765],seed[1963],seed[2234],seed[3483],seed[3492],seed[1181],seed[2040],seed[693],seed[3663],seed[3226],seed[80],seed[3858],seed[2783],seed[1723],seed[1309],seed[2834],seed[288],seed[1446],seed[673],seed[692],seed[524],seed[1808],seed[31],seed[2907],seed[3685],seed[1939],seed[3643],seed[262],seed[1087],seed[1173],seed[1191],seed[390],seed[3579],seed[2088],seed[2559],seed[2571],seed[2368],seed[3559],seed[1666],seed[771],seed[159],seed[686],seed[3340],seed[2803],seed[237],seed[474],seed[375],seed[1298],seed[1345],seed[3165],seed[2586],seed[2614],seed[117],seed[640],seed[3852],seed[1977],seed[3961],seed[68],seed[2513],seed[1978],seed[2310],seed[3211],seed[1097],seed[3997],seed[1217],seed[1900],seed[3304],seed[1731],seed[3728],seed[3332],seed[1449],seed[3703],seed[2157],seed[3975],seed[2014],seed[855],seed[191],seed[2983],seed[538],seed[817],seed[925],seed[2456],seed[1761],seed[2076],seed[839],seed[408],seed[3900],seed[1877],seed[984],seed[2546],seed[317],seed[3590],seed[2463],seed[2630],seed[1514],seed[3793],seed[2987],seed[949],seed[3956],seed[1659],seed[2300],seed[1709],seed[3693],seed[4059],seed[3880],seed[3248],seed[590],seed[2224],seed[749],seed[2148],seed[2609],seed[1581],seed[1973],seed[3071],seed[2991],seed[254],seed[550],seed[2284],seed[1494],seed[3690],seed[3555],seed[3792],seed[151],seed[661],seed[7],seed[2065],seed[4079],seed[2285],seed[89],seed[2740],seed[1760],seed[2664],seed[3051],seed[1568],seed[2489],seed[980],seed[2668],seed[1231],seed[1064],seed[3100],seed[3420],seed[3701],seed[236],seed[2728],seed[3901],seed[1347],seed[829],seed[3708],seed[2936],seed[3681],seed[3050],seed[2016],seed[754],seed[3996],seed[1924],seed[1935],seed[2169],seed[2925],seed[2106],seed[1754],seed[1705],seed[36],seed[3286],seed[115],seed[3625],seed[2336],seed[3292],seed[583],seed[713],seed[3206],seed[504],seed[603],seed[1743],seed[2391],seed[716],seed[2074],seed[1052],seed[2642],seed[3289],seed[3932],seed[3757],seed[2349],seed[1470],seed[3577],seed[2606],seed[4060],seed[3351],seed[3635],seed[709],seed[906],seed[2051],seed[3864],seed[3750],seed[3088],seed[152],seed[413],seed[1832],seed[894],seed[93],seed[2294],seed[3982],seed[1746],seed[1442],seed[2165],seed[3457],seed[3117],seed[823],seed[495],seed[1290],seed[2611],seed[2946],seed[2063],seed[3374],seed[2311],seed[427],seed[4036],seed[2205],seed[3946],seed[833],seed[1080],seed[2101],seed[3918],seed[475],seed[3496],seed[3473],seed[2078],seed[3250],seed[2382],seed[2090],seed[1511],seed[3623],seed[2100],seed[1382],seed[1966],seed[1437],seed[3922],seed[221],seed[122],seed[3732],seed[207],seed[4025],seed[3468],seed[1643],seed[2600],seed[3438],seed[2236],seed[653],seed[2568],seed[629],seed[1645],seed[2501],seed[1592],seed[2426],seed[601],seed[2174],seed[3834],seed[3525],seed[3278],seed[2757],seed[1482],seed[4054],seed[2721],seed[1342],seed[2251],seed[3556],seed[1458],seed[515],seed[2289],seed[1316],seed[931],seed[3613],seed[4094],seed[1928],seed[3879],seed[362],seed[767],seed[962],seed[882],seed[3515],seed[979],seed[2242],seed[2968],seed[71],seed[1364],seed[3821],seed[222],seed[844],seed[2510],seed[619],seed[1264],seed[537],seed[1938],seed[1265],seed[3406],seed[3794],seed[3427],seed[867],seed[1388],seed[2880],seed[513],seed[1344],seed[101],seed[1699],seed[69],seed[3333],seed[1407],seed[3935],seed[2001],seed[891],seed[3808],seed[4],seed[3674],seed[1542],seed[1902],seed[3948],seed[3352],seed[548],seed[233],seed[1679],seed[3315],seed[2635],seed[1378],seed[1190],seed[1013],seed[2226],seed[1668],seed[2842],seed[2974],seed[3077],seed[3495],seed[3986],seed[419],seed[3334],seed[3401],seed[1367],seed[3044],seed[2248],seed[1946],seed[585],seed[231],seed[1934],seed[1001],seed[1944],seed[169],seed[3570],seed[1138],seed[4045],seed[3419],seed[3228],seed[176],seed[2476],seed[3796],seed[617],seed[2469],seed[4068],seed[1234],seed[2542],seed[257],seed[2494],seed[3898],seed[2108],seed[3756],seed[1634],seed[1121],seed[3297],seed[2142],seed[2813],seed[3062],seed[1861],seed[1238],seed[274],seed[1164],seed[2158],seed[879],seed[3806],seed[976],seed[3797],seed[2839],seed[125],seed[1040],seed[3321],seed[3785],seed[3012],seed[3251],seed[2341],seed[3508],seed[706],seed[3549],seed[2785],seed[2605],seed[3507],seed[1045],seed[1120],seed[1755],seed[1600],seed[3715],seed[22],seed[1431],seed[828],seed[3589],seed[945],seed[211],seed[2824],seed[1764],seed[1654],seed[3480],seed[1226],seed[2570],seed[383],seed[1800],seed[2387],seed[1895],seed[761],seed[613],seed[3113],seed[1546],seed[3593],seed[1766],seed[311],seed[3096],seed[2821],seed[1871],seed[15],seed[973],seed[340],seed[3447],seed[3223],seed[2337],seed[734],seed[1018],seed[104],seed[3680],seed[1728],seed[3650],seed[3609],seed[3889],seed[3070],seed[2908],seed[2134],seed[303],seed[2191],seed[1621],seed[308],seed[747],seed[177],seed[996],seed[4014],seed[3531],seed[2487],seed[1438],seed[3778],seed[1562],seed[3087],seed[1884],seed[1420],seed[3911],seed[44],seed[2262],seed[3487],seed[974],seed[3436],seed[975],seed[2554],seed[249],seed[3709],seed[201],seed[553],seed[2374],seed[141],seed[2872],seed[3881],seed[1113],seed[267],seed[389],seed[2211],seed[1947],seed[2823],seed[1062],seed[2719],seed[2971],seed[1597],seed[2008],seed[1496],seed[3675],seed[845],seed[1330],seed[2859],seed[188],seed[1195],seed[195],seed[2539],seed[2961],seed[2046],seed[2155],seed[2825],seed[3482],seed[801],seed[57],seed[2215],seed[2527],seed[670],seed[4075],seed[3073],seed[1777],seed[3122],seed[2703],seed[50],seed[444],seed[3037],seed[663],seed[2905],seed[3859],seed[705],seed[2932],seed[2186],seed[3657],seed[372],seed[302],seed[874],seed[3943],seed[1220],seed[2117],seed[2563],seed[2738],seed[1157],seed[959],seed[624],seed[1397],seed[1452],seed[438],seed[3764],seed[508],seed[1368],seed[3963],seed[3239],seed[2071],seed[3772],seed[3469],seed[2124],seed[447],seed[2059],seed[1748],seed[1004],seed[24],seed[3150],seed[3448],seed[1910],seed[3972],seed[4021],seed[326],seed[840],seed[3153],seed[2895],seed[1839],seed[3342],seed[536],seed[2013],seed[227],seed[1396],seed[333],seed[501],seed[1661],seed[1433],seed[1375],seed[774],seed[3869],seed[2473],seed[98],seed[2295],seed[1209],seed[2449],seed[2268],seed[3256],seed[1398],seed[3345],seed[3554],seed[3103],seed[3714],seed[3390],seed[2389],seed[2095],seed[981],seed[3913],seed[2774],seed[3450],seed[4078],seed[234],seed[1208],seed[896],seed[493],seed[787],seed[4023],seed[3776],seed[162],seed[1094],seed[3843],seed[4027],seed[2885],seed[3947],seed[2362],seed[939],seed[2634],seed[2760],seed[3196],seed[445],seed[2779],seed[3568],seed[3016],seed[2753],seed[3544],seed[1314],seed[470],seed[2140],seed[3372],seed[3617],seed[3744],seed[2940],seed[531],seed[3017],seed[3743],seed[3446],seed[506],seed[2822],seed[3741],seed[1140],seed[872],seed[1640],seed[2712],seed[171],seed[2344],seed[3896],seed[837],seed[2988],seed[586],seed[2975],seed[2480],seed[12],seed[1472],seed[3300],seed[3824],seed[2394],seed[1451],seed[2316],seed[476],seed[2072],seed[731],seed[2596],seed[2705],seed[1631],seed[3275],seed[1851],seed[4064],seed[2044],seed[2937],seed[1782],seed[2835],seed[2941],seed[1214],seed[543],seed[3654],seed[2502],seed[1736],seed[1279],seed[2744],seed[750],seed[3973],seed[682],seed[3798],seed[2187],seed[1162],seed[446],seed[3031],seed[3414],seed[2432],seed[276],seed[414],seed[59],seed[206],seed[3486],seed[2963],seed[1642],seed[2271],seed[1333],seed[1948],seed[26],seed[730],seed[1797],seed[304],seed[1440],seed[23],seed[3089],seed[1971],seed[3546],seed[3355],seed[259],seed[450],seed[1727],seed[1584],seed[2496],seed[2581],seed[1655],seed[1297],seed[1422],seed[2620],seed[909],seed[3272],seed[2025],seed[18],seed[2276],seed[2659],seed[35],seed[741],seed[2641],seed[2281],seed[2317],seed[2686],seed[3160],seed[2010],seed[3039],seed[3320],seed[1512],seed[498],seed[161],seed[135],seed[1213],seed[2918],seed[1768],seed[782],seed[3652],seed[500],seed[2787],seed[789],seed[1391],seed[1036],seed[418],seed[3475],seed[2474],seed[755],seed[1586],seed[849],seed[2280],seed[3713],seed[205],seed[1188],seed[3676],seed[812],seed[1667],seed[2466],seed[2484],seed[834],seed[3576],seed[1613],seed[3435],seed[2221],seed[2578],seed[2452],seed[1976],seed[3207],seed[2229],seed[1685],seed[3527],seed[255],seed[2246],seed[1263],seed[433],seed[1007],seed[156],seed[598],seed[3519],seed[1002],seed[3758],seed[1756],seed[2379],seed[119],seed[2768],seed[2818],seed[1969],seed[1350],seed[3220],seed[2776],seed[1733],seed[2871],seed[2583],seed[1360],seed[1534],seed[3937],seed[407],seed[3698],seed[3354],seed[1530],seed[2650],seed[2655],seed[2329],seed[2624],seed[3586],seed[1975],seed[4081],seed[2325],seed[3179],seed[1480],seed[1960],seed[530],seed[2793],seed[2053],seed[223],seed[2862],seed[1583],seed[384],seed[2567],seed[79],seed[2942],seed[2837],seed[596],seed[429],seed[3873],seed[355],seed[1357],seed[2069],seed[929],seed[2367],seed[3751],seed[3430],seed[111],seed[1868],seed[490],seed[542],seed[3520],seed[780],seed[558],seed[3453],seed[1423],seed[2621],seed[2055],seed[3288],seed[2260],seed[2745],seed[3183],seed[1786],seed[1563],seed[2267],seed[3175],seed[2366],seed[1178],seed[3084],seed[1176],seed[3091],seed[3567],seed[1735],seed[668],seed[3979],seed[1092],seed[3021],seed[3296],seed[3841],seed[2841],seed[2577],seed[3455],seed[1750],seed[275],seed[3769],seed[3356],seed[2388],seed[3803],seed[1076],seed[3723],seed[189],seed[3561],seed[2402],seed[1379],seed[1504],seed[2881],seed[1880],seed[3886],seed[3056],seed[2322],seed[1793],seed[2675],seed[3945],seed[1617],seed[2427],seed[3988],seed[1171],seed[3734],seed[3162],seed[309],seed[271],seed[1386],seed[3009],seed[2509],seed[3648],seed[1381],seed[2067],seed[3558],seed[2081],seed[1089],seed[1010],seed[3121],seed[3562],seed[277],seed[282],seed[773],seed[1317],seed[3030],seed[1579],seed[435],seed[1558],seed[1827],seed[116],seed[963],seed[443],seed[1547],seed[3575],seed[1365],seed[2811],seed[1576],seed[1387],seed[2358],seed[647],seed[2365],seed[2762],seed[941],seed[3633],seed[426],seed[804],seed[2565],seed[1467],seed[3987],seed[3359],seed[2189],seed[1552],seed[3876],seed[3274],seed[948],seed[331],seed[3400],seed[480],seed[3209],seed[120],seed[2734],seed[2286],seed[252],seed[3266],seed[1858],seed[1812],seed[1455],seed[2461],seed[2731],seed[1032],seed[154],seed[656],seed[39],seed[3200],seed[202],seed[987],seed[1762],seed[337],seed[3086],seed[2663],seed[2769],seed[1463],seed[194],seed[3543],seed[886],seed[707],seed[1806],seed[3704],seed[2561],seed[82],seed[1838],seed[2162],seed[1477],seed[411],seed[3391],seed[784],seed[3441],seed[1759],seed[2984],seed[1326],seed[2043],seed[1184],seed[1956],seed[1593],seed[3168],seed[1261],seed[911],seed[1042],seed[283],seed[3669],seed[1869],seed[321],seed[3023],seed[134],seed[4086],seed[724],seed[2483],seed[1588],seed[552],seed[1564],seed[358],seed[2876],seed[1525],seed[2185],seed[198],seed[951],seed[2748],seed[600],seed[992],seed[3844],seed[2520],seed[1828],seed[1222],seed[1722],seed[1652],seed[3658],seed[2112],seed[606],seed[3962],seed[3809],seed[569],seed[1988],seed[3394],seed[1322],seed[3991],seed[792],seed[3404],seed[2220],seed[3388],seed[3638],seed[266],seed[109],seed[2278],seed[2352],seed[635],seed[3006],seed[224],seed[1738],seed[2377],seed[1696],seed[3326],seed[1307],seed[2345],seed[502],seed[1893],seed[3109],seed[2447],seed[347],seed[2493],seed[3688],seed[3025],seed[1732],seed[3361],seed[1675],seed[2441],seed[1879],seed[1225],seed[587],seed[1054],seed[208],seed[105],seed[463],seed[3152],seed[1840],seed[2350],seed[1193],seed[2660],seed[1487],seed[1392],seed[3072],seed[1686],seed[1949],seed[2315],seed[1131],seed[106],seed[76],seed[3959],seed[1159],seed[325],seed[1211],seed[3443],seed[3425],seed[2977],seed[2370],seed[2414],seed[299],seed[1249],seed[1836],seed[802],seed[166],seed[2404],seed[1077],seed[2674],seed[1351],seed[4090],seed[639],seed[1767],seed[1192],seed[577],seed[1031],seed[3246],seed[442],seed[559],seed[2622],seed[1158],seed[3260],seed[846],seed[863],seed[2764],seed[2526],seed[3382],seed[800],seed[1170],seed[3284],seed[2697],seed[3104],seed[3137],seed[1922],seed[1739],seed[1610],seed[2845],seed[2970],seed[2037],seed[146],seed[968],seed[3917],seed[1369],seed[3883],seed[2096],seed[3707],seed[2061],seed[3265],seed[3925],seed[3984],seed[1028],seed[4000],seed[58],seed[2020],seed[964],seed[1],seed[2116],seed[319],seed[1165],seed[671],seed[2792],seed[49],seed[1147],seed[4016],seed[1497],seed[952],seed[2595],seed[2193],seed[3594],seed[3990],seed[2123],seed[2153],seed[3258],seed[3412],seed[1468],seed[1641],seed[1522],seed[2864],seed[2160],seed[3370],seed[1997],seed[1473],seed[3465],seed[859],seed[1937],seed[2691],seed[2070],seed[320],seed[2105],seed[2816],seed[124],seed[999],seed[72],seed[3823],seed[612],seed[2425],seed[3142],seed[380],seed[1023],seed[1803],seed[3481],seed[534],seed[365],seed[2029],seed[1447],seed[901],seed[3636],seed[1638],seed[2506],seed[1503],seed[914],seed[3971],seed[17],seed[1874],seed[631],seed[514],seed[3934],seed[690],seed[4055],seed[2202],seed[338],seed[1908],seed[1204],seed[2766],seed[573],seed[2355],seed[1118],seed[3770],seed[1629],seed[842],seed[2591],seed[608],seed[2419],seed[3437],seed[1371],seed[1418],seed[334],seed[3134],seed[1289],seed[2802],seed[644],seed[3112],seed[3479],seed[1393],seed[1644],seed[1896],seed[1245],seed[938],seed[1243],seed[1259],seed[764],seed[1972],seed[3790],seed[1532],seed[2232],seed[597],seed[3369],seed[3565],seed[1246],seed[393],seed[3338],seed[3595],seed[1321],seed[8],seed[496],seed[2092],seed[648],seed[3392],seed[1704],seed[3553],seed[808],seed[1374],seed[3489],seed[3166],seed[1400],seed[3661],seed[2999],seed[1776],seed[3302],seed[1940],seed[243],seed[2312],seed[2739],seed[1936],seed[2245],seed[2024],seed[398],seed[1918],seed[2393],seed[4057],seed[1311],seed[505],seed[1366],seed[123],seed[3099],seed[3813],seed[770],seed[2515],seed[1421],seed[816],seed[2428],seed[2429],seed[4011],seed[3835],seed[2623],seed[431],seed[3736],seed[242],seed[2346],seed[3405],seed[3377],seed[4076],seed[1432],seed[565],seed[3171],seed[2168],seed[1135],seed[425],seed[1974],seed[3929],seed[1986],seed[2110],seed[4001],seed[3624],seed[2716],seed[1086],seed[3903],seed[3385],seed[1981],seed[3348],seed[1792],seed[1959],seed[4061],seed[1541],seed[1904],seed[432],seed[1656],seed[296],seed[1498],seed[291],seed[507],seed[2199],seed[462],seed[3994],seed[3645],seed[4041],seed[3472],seed[2726],seed[1464],seed[1660],seed[402],seed[1890],seed[3234],seed[2437],seed[184],seed[4092],seed[3204],seed[3173],seed[2438],seed[3902],seed[953],seed[2795],seed[424],seed[295],seed[1119],seed[2898],seed[2431],seed[638],seed[1276],seed[394],seed[3596],seed[2314],seed[461],seed[3832],seed[1932],seed[3862],seed[1434],seed[3389],seed[3235],seed[2514],seed[3920],seed[2633],seed[403],seed[3640],seed[1230],seed[1281],seed[1570],seed[676],seed[2254],seed[3213],seed[1107],seed[3422],seed[2482],seed[2299],seed[3182],seed[982],seed[2066],seed[1310],seed[575],seed[3860],seed[99],seed[95],seed[766],seed[3666],seed[1339],seed[1707],seed[621],seed[990],seed[1206],seed[858],seed[3060],seed[4088],seed[1987],seed[830],seed[2607],seed[2027],seed[777],seed[157],seed[1804],seed[4091],seed[1943],seed[3861],seed[636],seed[2498],seed[1299],seed[2866],seed[448],seed[2133],seed[3818],seed[3634],seed[1053],seed[248],seed[643],seed[102],seed[2773],seed[3067],seed[330],seed[3747],seed[4024],seed[2217],seed[2959],seed[1855],seed[1845],seed[1308],seed[56],seed[3146],seed[3667],seed[3916],seed[1110],seed[2952],seed[3999],seed[3605],seed[1239],seed[2518],seed[4043],seed[1809],seed[3777],seed[869],seed[391],seed[3444],seed[723],seed[1233],seed[1752],seed[2833],seed[3964],seed[2213],seed[270],seed[1484],seed[2468],seed[3215],seed[633],seed[2265],seed[2411],seed[3341],seed[457],seed[318],seed[3897],seed[936],seed[2877],seed[1215],seed[113],seed[3588],seed[2409],seed[2032],seed[3327],seed[881],seed[88],seed[192],seed[2640],seed[809],seed[3219],seed[250],seed[409],seed[1483],seed[3363],seed[1967],seed[3010],seed[3610],seed[153],seed[3057],seed[3157],seed[0],seed[342],seed[1267],seed[4071],seed[1538],seed[2424],seed[1508],seed[183],seed[2537],seed[3763],seed[2645],seed[428],seed[2207],seed[2588],seed[732],seed[3632],seed[3953],seed[3560],seed[3682],seed[2829],seed[185],seed[2852],seed[579],seed[3499],seed[1663],seed[720],seed[2395],seed[353],seed[287],seed[532],seed[2993],seed[694],seed[1030],seed[2652],seed[3819],seed[42],seed[3464],seed[813],seed[1533],seed[856],seed[2347],seed[3149],seed[1636],seed[3890],seed[306],seed[1907],seed[3306],seed[2843],seed[958],seed[3557],seed[2598],seed[1820],seed[3241],seed[1182],seed[5],seed[3653],seed[2684],seed[3622],seed[3116],seed[3221],seed[2896],seed[164],seed[1074],seed[1462],seed[3952],seed[3524],seed[832],seed[3339],seed[3915],seed[3065],seed[3598],seed[1850],seed[209],seed[3493],seed[3733],seed[1531],seed[3490],seed[1942],seed[2564],seed[2132],seed[1055],seed[3145],seed[2638],seed[3716],seed[3928]}),
        .cross_prob(cross_prob),
        .codeword(codeword12),
        .received(received12)
        );
    
    bsc bsc13(
        .clk(clk),
        .reset(reset),
        .seed({seed[2637],seed[694],seed[2721],seed[1265],seed[897],seed[3680],seed[2571],seed[1233],seed[866],seed[2447],seed[803],seed[536],seed[57],seed[827],seed[2742],seed[523],seed[305],seed[570],seed[1018],seed[33],seed[3448],seed[2408],seed[3419],seed[2792],seed[1566],seed[3413],seed[2068],seed[2167],seed[3122],seed[89],seed[1780],seed[1413],seed[3092],seed[858],seed[308],seed[2482],seed[2281],seed[2863],seed[251],seed[898],seed[855],seed[3575],seed[3080],seed[4023],seed[1322],seed[741],seed[149],seed[1258],seed[3555],seed[1677],seed[3383],seed[1578],seed[109],seed[3427],seed[1110],seed[2357],seed[239],seed[713],seed[3095],seed[309],seed[3628],seed[3664],seed[126],seed[379],seed[3140],seed[488],seed[1101],seed[3785],seed[3458],seed[3958],seed[3989],seed[2030],seed[3042],seed[103],seed[4020],seed[2595],seed[2188],seed[3604],seed[3607],seed[875],seed[2553],seed[1608],seed[260],seed[2183],seed[950],seed[1921],seed[359],seed[2265],seed[1557],seed[4039],seed[3154],seed[1231],seed[512],seed[2536],seed[147],seed[2170],seed[1889],seed[516],seed[2638],seed[915],seed[3250],seed[2052],seed[3356],seed[1073],seed[1562],seed[290],seed[3199],seed[2951],seed[2813],seed[2234],seed[1023],seed[3850],seed[3967],seed[3622],seed[3769],seed[697],seed[4043],seed[1296],seed[417],seed[1940],seed[792],seed[925],seed[3933],seed[1280],seed[2652],seed[276],seed[30],seed[2712],seed[2324],seed[3647],seed[3759],seed[3614],seed[1996],seed[3090],seed[1831],seed[2847],seed[1518],seed[1901],seed[2387],seed[2572],seed[3013],seed[2381],seed[2202],seed[2463],seed[157],seed[1136],seed[3948],seed[3873],seed[477],seed[2123],seed[232],seed[3313],seed[1631],seed[475],seed[1877],seed[1567],seed[1602],seed[1383],seed[2380],seed[220],seed[1686],seed[3502],seed[733],seed[1094],seed[2618],seed[2621],seed[3843],seed[775],seed[2740],seed[224],seed[2057],seed[3914],seed[375],seed[3959],seed[1708],seed[701],seed[911],seed[1180],seed[2133],seed[1038],seed[2418],seed[762],seed[1203],seed[1142],seed[2967],seed[254],seed[1432],seed[778],seed[1597],seed[568],seed[3477],seed[1282],seed[3827],seed[3161],seed[761],seed[184],seed[72],seed[228],seed[3976],seed[2020],seed[2707],seed[1556],seed[1834],seed[1174],seed[323],seed[98],seed[3182],seed[1781],seed[2877],seed[2431],seed[1320],seed[1793],seed[1181],seed[708],seed[1718],seed[1055],seed[3855],seed[2891],seed[3786],seed[441],seed[3815],seed[1267],seed[3936],seed[1473],seed[883],seed[2942],seed[2780],seed[4007],seed[1712],seed[3611],seed[1930],seed[2100],seed[3789],seed[3469],seed[1040],seed[2991],seed[3816],seed[2968],seed[1157],seed[1255],seed[979],seed[362],seed[110],seed[3739],seed[1010],seed[3303],seed[2625],seed[2474],seed[2770],seed[91],seed[2285],seed[3861],seed[3610],seed[3943],seed[1974],seed[3990],seed[1873],seed[661],seed[1008],seed[2500],seed[3652],seed[3937],seed[1962],seed[1495],seed[455],seed[1199],seed[2749],seed[2522],seed[2062],seed[1498],seed[3633],seed[1421],seed[2042],seed[2870],seed[2289],seed[2101],seed[3973],seed[3545],seed[798],seed[1293],seed[1559],seed[142],seed[1049],seed[2376],seed[404],seed[3314],seed[1388],seed[3075],seed[206],seed[1735],seed[3218],seed[3508],seed[3475],seed[2636],seed[3297],seed[526],seed[2475],seed[1170],seed[2941],seed[2731],seed[3594],seed[2643],seed[394],seed[1749],seed[696],seed[751],seed[3236],seed[3845],seed[2850],seed[2450],seed[4022],seed[2581],seed[1381],seed[1342],seed[2110],seed[175],seed[583],seed[808],seed[3134],seed[2327],seed[581],seed[3162],seed[2527],seed[3022],seed[6],seed[3331],seed[918],seed[3821],seed[1980],seed[3187],seed[2868],seed[386],seed[2141],seed[1493],seed[3328],seed[1818],seed[1364],seed[3893],seed[2488],seed[2258],seed[569],seed[1088],seed[2006],seed[2921],seed[3569],seed[557],seed[2095],seed[1738],seed[1347],seed[1403],seed[1987],seed[73],seed[1273],seed[3320],seed[2341],seed[2524],seed[3995],seed[3773],seed[69],seed[2270],seed[1279],seed[47],seed[2650],seed[90],seed[1451],seed[3077],seed[3979],seed[2689],seed[2913],seed[233],seed[2660],seed[182],seed[2144],seed[1066],seed[2119],seed[85],seed[92],seed[1097],seed[3412],seed[1439],seed[2084],seed[3846],seed[594],seed[3694],seed[108],seed[3919],seed[2980],seed[2125],seed[3315],seed[511],seed[1852],seed[352],seed[1392],seed[1540],seed[447],seed[3798],seed[3033],seed[1804],seed[2701],seed[61],seed[3782],seed[3517],seed[1574],seed[2292],seed[2129],seed[3145],seed[2746],seed[1747],seed[3925],seed[2287],seed[650],seed[1569],seed[2237],seed[2348],seed[373],seed[2074],seed[2458],seed[3568],seed[1946],seed[1515],seed[3209],seed[2692],seed[3668],seed[1299],seed[1437],seed[2817],seed[1806],seed[784],seed[498],seed[3757],seed[1648],seed[1820],seed[1630],seed[2412],seed[2319],seed[3868],seed[102],seed[508],seed[2768],seed[363],seed[3358],seed[3533],seed[912],seed[1799],seed[158],seed[2139],seed[3091],seed[3118],seed[873],seed[481],seed[29],seed[2539],seed[1212],seed[2986],seed[1918],seed[1898],seed[3345],seed[112],seed[3999],seed[2670],seed[948],seed[1828],seed[3335],seed[4008],seed[3509],seed[3360],seed[2704],seed[3440],seed[1645],seed[3120],seed[3932],seed[118],seed[757],seed[1797],seed[2711],seed[2104],seed[2714],seed[3210],seed[3205],seed[3025],seed[2912],seed[1007],seed[1655],seed[3691],seed[3586],seed[974],seed[3649],seed[1813],seed[544],seed[1976],seed[3423],seed[3188],seed[2212],seed[3211],seed[470],seed[3044],seed[1414],seed[3825],seed[947],seed[2346],seed[1458],seed[861],seed[1048],seed[3808],seed[2487],seed[848],seed[1098],seed[3130],seed[2051],seed[3975],seed[530],seed[1394],seed[2282],seed[3168],seed[1145],seed[3981],seed[2184],seed[2111],seed[395],seed[1395],seed[1721],seed[646],seed[2145],seed[351],seed[760],seed[2448],seed[2804],seed[3651],seed[237],seed[3201],seed[2113],seed[3666],seed[2869],seed[563],seed[2047],seed[3253],seed[288],seed[4001],seed[3867],seed[2254],seed[3641],seed[2858],seed[2932],seed[2723],seed[155],seed[2117],seed[41],seed[3831],seed[3325],seed[3333],seed[2922],seed[3219],seed[871],seed[1298],seed[1295],seed[2286],seed[1512],seed[2601],seed[3112],seed[83],seed[407],seed[1489],seed[2955],seed[1922],seed[944],seed[2541],seed[1288],seed[3105],seed[2271],seed[1917],seed[125],seed[1585],seed[3116],seed[2089],seed[1639],seed[2401],seed[3707],seed[2881],seed[926],seed[689],seed[3059],seed[436],seed[1925],seed[1244],seed[2058],seed[1990],seed[1125],seed[494],seed[2432],seed[4015],seed[1727],seed[3903],seed[1459],seed[1270],seed[3896],seed[2681],seed[2493],seed[1874],seed[1152],seed[657],seed[1189],seed[774],seed[221],seed[88],seed[3506],seed[3587],seed[200],seed[3483],seed[3035],seed[3371],seed[723],seed[3336],seed[1767],seed[905],seed[2366],seed[1651],seed[1341],seed[981],seed[2895],seed[1324],seed[687],seed[458],seed[3904],seed[2873],seed[1812],seed[3444],seed[3365],seed[921],seed[1571],seed[3052],seed[3408],seed[844],seed[319],seed[946],seed[3257],seed[3326],seed[1359],seed[1993],seed[2176],seed[2229],seed[2027],seed[3576],seed[1503],seed[2739],seed[1609],seed[2166],seed[3573],seed[2120],seed[2186],seed[261],seed[2717],seed[1740],seed[623],seed[1337],seed[2733],seed[339],seed[3504],seed[52],seed[2853],seed[3269],seed[1915],seed[3623],seed[3179],seed[1287],seed[4049],seed[3447],seed[3196],seed[549],seed[1286],seed[1128],seed[3086],seed[2426],seed[2677],seed[2501],seed[195],seed[2140],seed[3180],seed[1967],seed[1722],seed[1241],seed[879],seed[919],seed[1884],seed[1448],seed[1348],seed[3501],seed[138],seed[3947],seed[1516],seed[3629],seed[2776],seed[585],seed[3830],seed[695],seed[1688],seed[1961],seed[1469],seed[1294],seed[3701],seed[3688],seed[78],seed[3912],seed[137],seed[1719],seed[3512],seed[4014],seed[1254],seed[2800],seed[2886],seed[2259],seed[489],seed[2180],seed[2971],seed[2159],seed[2230],seed[1452],seed[3980],seed[2889],seed[3050],seed[3390],seed[2726],seed[66],seed[425],seed[133],seed[3388],seed[3391],seed[296],seed[3363],seed[3318],seed[727],seed[3164],seed[1785],seed[2112],seed[3375],seed[3535],seed[1202],seed[2196],seed[1616],seed[3171],seed[304],seed[1981],seed[3456],seed[3340],seed[439],seed[3415],seed[122],seed[3245],seed[1568],seed[3418],seed[360],seed[2065],seed[3730],seed[1118],seed[3395],seed[1752],seed[4086],seed[2861],seed[2149],seed[1166],seed[1120],seed[1851],seed[344],seed[592],seed[1580],seed[2339],seed[4012],seed[824],seed[3378],seed[144],seed[3791],seed[3818],seed[2856],seed[3264],seed[2702],seed[1237],seed[924],seed[2328],seed[1307],seed[2969],seed[1302],seed[2729],seed[53],seed[2246],seed[2538],seed[2419],seed[1988],seed[3767],seed[1809],seed[752],seed[3494],seed[1496],seed[411],seed[3076],seed[160],seed[1283],seed[2513],seed[940],seed[2175],seed[3765],seed[3716],seed[3638],seed[3267],seed[445],seed[95],seed[2083],seed[434],seed[448],seed[586],seed[3918],seed[1937],seed[1031],seed[759],seed[2152],seed[2477],seed[2273],seed[1576],seed[1702],seed[747],seed[2178],seed[719],seed[3811],seed[505],seed[665],seed[1973],seed[3372],seed[3015],seed[856],seed[1129],seed[484],seed[572],seed[2795],seed[3580],seed[2480],seed[2005],seed[3030],seed[2959],seed[2245],seed[1637],seed[259],seed[966],seed[3175],seed[1509],seed[2018],seed[2546],seed[3141],seed[982],seed[2761],seed[2405],seed[3554],seed[2478],seed[4072],seed[1099],seed[1113],seed[3528],seed[471],seed[1054],seed[2741],seed[3754],seed[2748],seed[1153],seed[3183],seed[1205],seed[3630],seed[3910],seed[2848],seed[870],seed[1778],seed[3747],seed[1084],seed[3496],seed[2250],seed[1319],seed[2266],seed[216],seed[1904],seed[1697],seed[2439],seed[3087],seed[2168],seed[1275],seed[2686],seed[4069],seed[1215],seed[217],seed[1433],seed[2845],seed[266],seed[653],seed[3146],seed[1707],seed[1162],seed[1005],seed[3834],seed[226],seed[630],seed[3058],seed[1528],seed[3272],seed[4077],seed[3480],seed[113],seed[2011],seed[2617],seed[3338],seed[3471],seed[4004],seed[1742],seed[3881],seed[189],seed[1179],seed[816],seed[1570],seed[1882],seed[4030],seed[3824],seed[1382],seed[3829],seed[2375],seed[1788],seed[1543],seed[3616],seed[1938],seed[614],seed[1680],seed[2841],seed[1713],seed[2197],seed[2545],seed[1530],seed[348],seed[4085],seed[2972],seed[2523],seed[989],seed[1687],seed[2658],seed[3278],seed[1832],seed[928],seed[3160],seed[3439],seed[26],seed[2404],seed[491],seed[3813],seed[1160],seed[3810],seed[1126],seed[4092],seed[4024],seed[1815],seed[2451],seed[185],seed[3273],seed[32],seed[2263],seed[2903],seed[3317],seed[2521],seed[401],seed[2803],seed[3312],seed[769],seed[2774],seed[2472],seed[4038],seed[3300],seed[2878],seed[1027],seed[4050],seed[1367],seed[2751],seed[3865],seed[190],seed[3887],seed[3069],seed[887],seed[3978],seed[3957],seed[952],seed[2081],seed[2876],seed[3485],seed[467],seed[3894],seed[954],seed[3064],seed[1720],seed[1075],seed[988],seed[515],seed[294],seed[2126],seed[63],seed[1711],seed[1067],seed[1971],seed[2824],seed[287],seed[1634],seed[1632],seed[1816],seed[3961],seed[616],seed[3492],seed[4010],seed[3942],seed[3531],seed[2198],seed[2283],seed[1551],seed[3909],seed[3429],seed[2135],seed[1186],seed[1600],seed[151],seed[2767],seed[1524],seed[3321],seed[3566],seed[1859],seed[3732],seed[3299],seed[909],seed[2840],seed[4047],seed[1610],seed[1964],seed[2732],seed[2516],seed[474],seed[524],seed[1091],seed[1340],seed[1256],seed[2703],seed[1150],seed[238],seed[793],seed[1879],seed[3343],seed[393],seed[114],seed[3561],seed[3579],seed[2849],seed[3449],seed[763],seed[1053],seed[4087],seed[1979],seed[148],seed[818],seed[3493],seed[2974],seed[1844],seed[1042],seed[613],seed[2148],seed[3734],seed[3750],seed[3593],seed[2954],seed[2326],seed[3702],seed[2651],seed[1857],seed[2679],seed[2910],seed[503],seed[256],seed[2044],seed[490],seed[2568],seed[100],seed[3800],seed[2189],seed[865],seed[3653],seed[183],seed[2818],seed[2136],seed[2305],seed[1044],seed[2407],seed[343],seed[1345],seed[50],seed[2243],seed[2709],seed[656],seed[3037],seed[2438],seed[336],seed[2543],seed[1374],seed[1969],seed[150],seed[1717],seed[3968],seed[3479],seed[746],seed[2783],seed[1855],seed[1537],seed[2471],seed[3753],seed[212],seed[850],seed[2037],seed[2008],seed[1449],seed[2616],seed[1856],seed[1491],seed[2436],seed[1285],seed[1513],seed[231],seed[755],seed[2984],seed[4091],seed[2570],seed[1725],seed[3807],seed[1849],seed[1590],seed[878],seed[2116],seed[3373],seed[3931],seed[1839],seed[1024],seed[3073],seed[3450],seed[2278],seed[2675],seed[671],seed[4074],seed[284],seed[1032],seed[3008],seed[3783],seed[2156],seed[1309],seed[560],seed[2316],seed[2187],seed[584],seed[1692],seed[3591],seed[198],seed[2288],seed[1396],seed[1850],seed[3403],seed[3525],seed[3115],seed[839],seed[2866],seed[428],seed[1245],seed[2452],seed[3156],seed[3268],seed[935],seed[19],seed[3900],seed[2384],seed[4002],seed[3776],seed[3292],seed[3377],seed[1490],seed[3930],seed[2620],seed[3128],seed[1953],seed[1910],seed[380],seed[3712],seed[2342],seed[1625],seed[3152],seed[649],seed[2907],seed[2276],seed[3203],seed[2661],seed[2730],seed[2309],seed[1483],seed[575],seed[3812],seed[2103],seed[3874],seed[3433],seed[501],seed[4036],seed[1249],seed[3571],seed[3287],seed[652],seed[76],seed[11],seed[2576],seed[3640],seed[3244],seed[1221],seed[1488],seed[1714],seed[3693],seed[2079],seed[662],seed[2077],seed[2397],seed[3157],seed[120],seed[2574],seed[2470],seed[4018],seed[84],seed[2777],seed[194],seed[1658],seed[1021],seed[1661],seed[1592],seed[1529],seed[3212],seed[885],seed[2865],seed[3728],seed[2540],seed[1045],seed[1681],seed[2585],seed[443],seed[4000],seed[2605],seed[2512],seed[3498],seed[3913],seed[209],seed[215],seed[2389],seed[3478],seed[2765],seed[922],seed[1734],seed[893],seed[163],seed[1071],seed[2495],seed[204],seed[459],seed[3537],seed[3663],seed[3240],seed[1028],seed[622],seed[3858],seed[3016],seed[3998],seed[3549],seed[2678],seed[1517],seed[2157],seed[4042],seed[881],seed[2925],seed[3070],seed[1754],seed[833],seed[1866],seed[3165],seed[749],seed[387],seed[3281],seed[642],seed[1497],seed[2952],seed[1876],seed[1875],seed[104],seed[3705],seed[250],seed[2093],seed[1934],seed[2799],seed[3768],seed[1078],seed[3167],seed[3715],seed[3801],seed[3627],seed[862],seed[3286],seed[2359],seed[1111],seed[1304],seed[4059],seed[1885],seed[1903],seed[3905],seed[107],seed[1694],seed[886],seed[3047],seed[2429],seed[976],seed[329],seed[2628],seed[2990],seed[3645],seed[680],seed[3302],seed[1746],seed[3686],seed[1363],seed[3305],seed[1741],seed[2199],seed[2299],seed[4057],seed[285],seed[242],seed[135],seed[2734],seed[2530],seed[1272],seed[2544],seed[2534],seed[2988],seed[3259],seed[1362],seed[1508],seed[1278],seed[2838],seed[1886],seed[3421],seed[1899],seed[1246],seed[1914],seed[1614],seed[2078],seed[2274],seed[2899],seed[12],seed[1739],seed[1002],seed[2242],seed[1191],seed[2191],seed[1243],seed[1116],seed[3396],seed[3382],seed[3],seed[2267],seed[1184],seed[2964],seed[229],seed[2607],seed[3949],seed[1108],seed[2713],seed[2331],seed[45],seed[2944],seed[3114],seed[3847],seed[998],seed[1888],seed[509],seed[571],seed[1554],seed[3578],seed[1823],seed[193],seed[1313],seed[1006],seed[1092],seed[235],seed[2473],seed[1536],seed[1138],seed[3654],seed[1555],seed[2798],seed[1628],seed[3956],seed[2094],seed[1505],seed[2115],seed[685],seed[2494],seed[2611],seed[202],seed[3915],seed[3232],seed[1761],seed[2771],seed[1972],seed[1195],seed[3696],seed[927],seed[3615],seed[2209],seed[655],seed[1955],seed[1081],seed[1864],seed[2306],seed[3697],seed[3362],seed[3608],seed[161],seed[2253],seed[3366],seed[1690],seed[2823],seed[2815],seed[754],seed[3417],seed[1957],seed[3039],seed[1247],seed[3227],seed[958],seed[1706],seed[3970],seed[3256],seed[543],seed[181],seed[3597],seed[1629],seed[2950],seed[3738],seed[620],seed[632],seed[410],seed[264],seed[3005],seed[821],seed[2039],seed[660],seed[2363],seed[500],seed[2185],seed[1626],seed[3246],seed[1748],seed[3006],seed[36],seed[553],seed[2846],seed[3529],seed[782],seed[2213],seed[1466],seed[2067],seed[3987],seed[1223],seed[96],seed[1709],seed[1698],seed[2926],seed[3177],seed[1956],seed[1867],seed[3637],seed[2710],seed[2313],seed[3584],seed[2232],seed[3612],seed[442],seed[3908],seed[369],seed[3662],seed[1519],seed[3119],seed[1950],seed[535],seed[2593],seed[3117],seed[1660],seed[3271],seed[2708],seed[3406],seed[1532],seed[3319],seed[1346],seed[1220],seed[3606],seed[2464],seed[2511],seed[3247],seed[74],seed[3195],seed[1595],seed[3658],seed[539],seed[1573],seed[3676],seed[403],seed[1970],seed[907],seed[3216],seed[2457],seed[366],seed[2296],seed[610],seed[809],seed[3027],seed[3735],seed[3720],seed[2097],seed[440],seed[3137],seed[3266],seed[1486],seed[1426],seed[2754],seed[328],seed[1482],seed[542],seed[1586],seed[1306],seed[1375],seed[1649],seed[3842],seed[2592],seed[580],seed[3283],seed[949],seed[303],seed[559],seed[3139],seed[2160],seed[3899],seed[2696],seed[2551],seed[178],seed[2904],seed[2936],seed[3742],seed[2307],seed[1531],seed[3285],seed[247],seed[2997],seed[2216],seed[3428],seed[293],seed[851],seed[3660],seed[2354],seed[2619],seed[1161],seed[3710],seed[2090],seed[3135],seed[3692],seed[3101],seed[838],seed[3397],seed[2608],seed[2982],seed[2021],seed[651],seed[3552],seed[2193],seed[628],seed[2315],seed[2531],seed[3648],seed[3558],seed[332],seed[771],seed[124],seed[270],seed[3675],seed[3851],seed[3771],seed[1881],seed[902],seed[1263],seed[2023],seed[546],seed[268],seed[2303],seed[2165],seed[2034],seed[3222],seed[207],seed[659],seed[277],seed[4065],seed[2872],seed[1615],seed[1906],seed[408],seed[2181],seed[3598],seed[1004],seed[1807],seed[3214],seed[146],seed[334],seed[959],seed[2888],seed[3011],seed[3826],seed[1544],seed[1526],seed[3426],seed[1100],seed[48],seed[1271],seed[2781],seed[418],seed[1774],seed[764],seed[188],seed[1646],seed[3174],seed[1253],seed[4066],seed[2340],seed[3736],seed[768],seed[3354],seed[2559],seed[2484],seed[2075],seed[2535],seed[1039],seed[548],seed[3169],seed[1082],seed[1547],seed[506],seed[4073],seed[3010],seed[3308],seed[492],seed[731],seed[1281],seed[1941],seed[337],seed[4089],seed[3155],seed[1926],seed[639],seed[22],seed[1389],seed[244],seed[996],seed[3526],seed[1998],seed[2409],seed[564],seed[1182],seed[132],seed[521],seed[2879],seed[307],seed[94],seed[1463],seed[3996],seed[888],seed[895],seed[1034],seed[3822],seed[3809],seed[3054],seed[116],seed[578],seed[3107],seed[4076],seed[579],seed[2312],seed[3237],seed[801],seed[396],seed[1290],seed[1035],seed[2355],seed[683],seed[1982],seed[1366],seed[811],seed[2134],seed[2802],seed[1456],seed[2343],seed[1619],seed[2885],seed[376],seed[3323],seed[1724],seed[3001],seed[2422],seed[2060],seed[1887],seed[3194],seed[1977],seed[2589],seed[111],seed[3066],seed[2639],seed[40],seed[3024],seed[3983],seed[3176],seed[3729],seed[3096],seed[3793],seed[3003],seed[1012],seed[2003],seed[1656],seed[34],seed[419],seed[2758],seed[1442],seed[2374],seed[1939],seed[882],seed[60],seed[3743],seed[2719],seed[2007],seed[1894],seed[3746],seed[3225],seed[599],seed[2421],seed[540],seed[27],seed[21],seed[3906],seed[3113],seed[3950],seed[829],seed[2855],seed[44],seed[278],seed[3724],seed[3596],seed[1783],seed[736],seed[3055],seed[2322],seed[514],seed[867],seed[1331],seed[3346],seed[3048],seed[1443],seed[1444],seed[169],seed[2364],seed[3466],seed[240],seed[3191],seed[3136],seed[1172],seed[3656],seed[1447],seed[1222],seed[3941],seed[1151],seed[3088],seed[3684],seed[2162],seed[3499],seed[814],seed[2820],seed[82],seed[799],seed[658],seed[3282],seed[3089],seed[1699],seed[2901],seed[2102],seed[1891],seed[2537],seed[997],seed[711],seed[758],seed[2793],seed[674],seed[370],seed[1905],seed[987],seed[1336],seed[1975],seed[218],seed[681],seed[4028],seed[3971],seed[1732],seed[3327],seed[1208],seed[438],seed[1323],seed[199],seed[1207],seed[3550],seed[2252],seed[3374],seed[720],seed[3885],seed[1214],seed[2498],seed[1771],seed[2467],seed[2843],seed[2909],seed[345],seed[2555],seed[3437],seed[1252],seed[3489],seed[3238],seed[2206],seed[4082],seed[1434],seed[4071],seed[3260],seed[537],seed[611],seed[1377],seed[3065],seed[1015],seed[2029],seed[2578],seed[1908],seed[3962],seed[3784],seed[4078],seed[3142],seed[2829],seed[1438],seed[3324],seed[2138],seed[706],seed[86],seed[2900],seed[3231],seed[1404],seed[1502],seed[702],seed[480],seed[1058],seed[2667],seed[3422],seed[2132],seed[1315],seed[3307],seed[1134],seed[3208],seed[1485],seed[1931],seed[971],seed[3491],seed[1504],seed[263],seed[1037],seed[2143],seed[2425],seed[1653],seed[1462],seed[2565],seed[3229],seed[3505],seed[3560],seed[3460],seed[1617],seed[325],seed[2688],seed[2588],seed[3543],seed[2241],seed[1096],seed[283],seed[2012],seed[728],seed[2264],seed[3452],seed[1830],seed[2054],seed[2778],seed[890],seed[2587],seed[2979],seed[3988],seed[51],seed[1117],seed[2836],seed[2646],seed[2987],seed[1399],seed[3602],seed[1301],seed[806],seed[3018],seed[2515],seed[3572],seed[740],seed[2382],seed[1772],seed[413],seed[3565],seed[3524],seed[364],seed[1511],seed[2875],seed[3751],seed[1932],seed[2594],seed[1453],seed[248],seed[615],seed[3657],seed[2529],seed[3060],seed[703],seed[357],seed[2573],seed[1072],seed[589],seed[1318],seed[174],seed[1642],seed[3643],seed[59],seed[3520],seed[3019],seed[1405],seed[2158],seed[469],seed[783],seed[933],seed[2017],seed[3454],seed[507],seed[551],seed[2221],seed[437],seed[555],seed[1520],seed[2000],seed[682],seed[1919],seed[3590],seed[2549],seed[2256],seed[2469],seed[2240],seed[2934],seed[3802],seed[2455],seed[4009],seed[1907],seed[2066],seed[4063],seed[291],seed[3953],seed[1095],seed[1327],seed[2064],seed[2235],seed[1836],seed[2417],seed[1123],seed[4090],seed[3002],seed[3848],seed[3974],seed[874],seed[286],seed[825],seed[3921],seed[1169],seed[3965],seed[1929],seed[2174],seed[2598],seed[3562],seed[2466],seed[2508],seed[734],seed[3511],seed[2718],seed[3659],seed[2687],seed[2414],seed[1696],seed[2356],seed[666],seed[3547],seed[2649],seed[3582],seed[1211],seed[637],seed[1542],seed[87],seed[3553],seed[3780],seed[518],seed[744],seed[1065],seed[2812],seed[1481],seed[127],seed[1158],seed[371],seed[3446],seed[1356],seed[3226],seed[1292],seed[1952],seed[3288],seed[392],seed[4095],seed[1057],seed[1784],seed[2153],seed[117],seed[3410],seed[3067],seed[300],seed[1026],seed[2244],seed[486],seed[1124],seed[2806],seed[1579],seed[1330],seed[3393],seed[3837],seed[3849],seed[612],seed[1693],seed[3760],seed[3669],seed[619],seed[4061],seed[1127],seed[1277],seed[1733],seed[2349],seed[2828],seed[3513],seed[820],seed[317],seed[576],seed[2410],seed[279],seed[1417],seed[3515],seed[2172],seed[1751],seed[3519],seed[341],seed[3166],seed[2514],seed[1763],seed[2070],seed[3839],seed[1352],seed[2373],seed[1043],seed[2350],seed[969],seed[208],seed[2706],seed[435],seed[3772],seed[3028],seed[3293],seed[2844],seed[3009],seed[2251],seed[698],seed[1627],seed[2906],seed[2599],seed[2096],seed[2329],seed[3451],seed[931],seed[16],seed[729],seed[673],seed[2561],seed[3261],seed[3945],seed[2837],seed[302],seed[957],seed[3880],seed[2519],seed[3476],seed[3852],seed[267],seed[2001],seed[1479],seed[1685],seed[213],seed[3193],seed[201],seed[3674],seed[1782],seed[1033],seed[2128],seed[1450],seed[3051],seed[1177],seed[2965],seed[3540],seed[4053],seed[1845],seed[1467],seed[1022],seed[454],seed[1548],seed[4068],seed[2632],seed[192],seed[2640],seed[1703],seed[3538],seed[795],seed[1052],seed[725],seed[3098],seed[1942],seed[18],seed[1726],seed[167],seed[2773],seed[942],seed[1470],seed[1471],seed[3392],seed[3523],seed[2489],seed[667],seed[2272],seed[910],seed[3764],seed[3626],seed[2736],seed[3123],seed[605],seed[1923],seed[2927],seed[863],seed[3866],seed[609],seed[3939],seed[2919],seed[269],seed[2295],seed[2669],seed[2291],seed[3275],seed[2962],seed[361],seed[3311],seed[1863],seed[1476],seed[2930],seed[2975],seed[624],seed[716],seed[1200],seed[2775],seed[776],seed[1606],seed[1549],seed[3559],seed[937],seed[2190],seed[2591],seed[3255],seed[3876],seed[787],seed[2961],seed[2600],seed[1912],seed[1730],seed[177],seed[2908],seed[1155],seed[627],seed[1076],seed[3097],seed[995],seed[3725],seed[1670],seed[1020],seed[281],seed[3796],seed[1563],seed[3964],seed[2437],seed[2918],seed[1840],seed[2610],seed[2154],seed[3721],seed[691],seed[1135],seed[1368],seed[608],seed[1829],seed[1985],seed[930],seed[2786],seed[1995],seed[3411],seed[1847],seed[2171],seed[714],seed[2108],seed[2393],seed[994],seed[1173],seed[934],seed[2635],seed[837],seed[153],seed[3886],seed[2146],seed[1525],seed[2105],seed[3871],seed[17],seed[3551],seed[289],seed[1872],seed[1425],seed[346],seed[4034],seed[3711],seed[1001],seed[3642],seed[3138],seed[1090],seed[1349],seed[2131],seed[1787],seed[1227],seed[826],seed[2],seed[2832],seed[4048],seed[3744],seed[3486],seed[3023],seed[3530],seed[3040],seed[450],seed[3034],seed[648],seed[4031],seed[1494],seed[2035],seed[4081],seed[3779],seed[1539],seed[3546],seed[943],seed[941],seed[128],seed[203],seed[2928],seed[3085],seed[1046],seed[872],seed[1700],seed[2896],seed[750],seed[3280],seed[25],seed[3698],seed[1657],seed[3198],seed[2043],seed[2092],seed[3963],seed[241],seed[2580],seed[2724],seed[415],seed[1361],seed[2998],seed[420],seed[960],seed[1080],seed[1623],seed[2978],seed[1933],seed[1289],seed[2905],seed[3589],seed[1800],seed[1764],seed[222],seed[565],seed[3761],seed[1682],seed[3683],seed[2563],seed[2280],seed[601],seed[2462],seed[3984],seed[186],seed[2575],seed[3386],seed[1947],seed[2835],seed[1596],seed[3790],seed[1750],seed[405],seed[721],seed[1613],seed[2630],seed[2400],seed[3817],seed[1790],seed[2890],seed[510],seed[381],seed[426],seed[1115],seed[3516],seed[1861],seed[2444],seed[3402],seed[678],seed[2238],seed[67],seed[3536],seed[1014],seed[1268],seed[3126],seed[2631],seed[3352],seed[3353],seed[1801],seed[2923],seed[173],seed[1047],seed[2325],seed[2031],seed[3869],seed[1621],seed[3057],seed[139],seed[39],seed[3290],seed[929],seed[1062],seed[1064],seed[2615],seed[3841],seed[2371],seed[2087],seed[903],seed[3111],seed[991],seed[2388],seed[3681],seed[2249],seed[37],seed[1167],seed[2973],seed[1593],seed[2490],seed[2048],seed[3541],seed[3709],seed[823],seed[301],seed[3084],seed[1779],seed[1729],seed[3892],seed[840],seed[1860],seed[0],seed[1365],seed[4021],seed[3110],seed[3158],seed[1089],seed[451],seed[1583],seed[457],seed[2874],seed[2779],seed[2173],seed[1997],seed[2526],seed[1197],seed[430],seed[1354],seed[65],seed[849],seed[3109],seed[1079],seed[3708],seed[3888],seed[93],seed[1016],seed[726],seed[1219],seed[1564],seed[1920],seed[2914],seed[3507],seed[965],seed[1407],seed[1674],seed[311],seed[2558],seed[1704],seed[2301],seed[2764],seed[115],seed[633],seed[2269],seed[3349],seed[4017],seed[1178],seed[1871],seed[1013],seed[1461],seed[1604],seed[3986],seed[3355],seed[2161],seed[3854],seed[3376],seed[3230],seed[3436],seed[236],seed[1063],seed[347],seed[917],seed[3603],seed[2690],seed[1140],seed[3459],seed[2468],seed[3241],seed[2496],seed[2685],seed[3472],seed[14],seed[1107],seed[868],seed[479],seed[3342],seed[2169],seed[1410],seed[906],seed[1441],seed[1499],seed[3197],seed[499],seed[1297],seed[28],seed[3689],seed[2333],seed[2697],seed[1343],seed[1011],seed[1507],seed[2217],seed[1880],seed[3254],seed[1500],seed[2377],seed[1652],seed[2107],seed[3178],seed[2787],seed[2204],seed[2528],seed[3733],seed[828],seed[2195],seed[3014],seed[1445],seed[1715],seed[900],seed[140],seed[1538],seed[2369],seed[3726],seed[2406],seed[2948],seed[3723],seed[1419],seed[3351],seed[836],seed[1546],seed[1335],seed[796],seed[834],seed[3857],seed[79],seed[2819],seed[449],seed[1984],seed[2737],seed[846],seed[1676],seed[3838],seed[669],seed[4005],seed[789],seed[901],seed[1777],seed[3994],seed[3737],seed[1131],seed[1429],seed[2399],seed[2441],seed[1316],seed[1753],seed[3079],seed[141],seed[1259],seed[1475],seed[522],seed[3316],seed[1406],seed[3190],seed[3542],seed[3289],seed[1662],seed[1228],seed[2810],seed[745],seed[832],seed[1059],seed[2569],seed[2360],seed[1669],seed[735],seed[629],seed[2378],seed[9],seed[590],seed[4019],seed[748],seed[1165],seed[3279],seed[3882],seed[2233],seed[3699],seed[3357],seed[3017],seed[3424],seed[2759],seed[62],seed[1112],seed[2634],seed[271],seed[3670],seed[1074],seed[772],seed[587],seed[2673],seed[2362],seed[986],seed[1792],seed[1386],seed[554],seed[797],seed[2834],seed[2791],seed[1185],seed[3159],seed[779],seed[472],seed[3147],seed[2808],seed[1594],seed[2228],seed[1892],seed[3094],seed[1527],seed[3510],seed[2150],seed[1262],seed[990],seed[1913],seed[3778],seed[2368],seed[1701],seed[3129],seed[4080],seed[4052],seed[1759],seed[282],seed[1371],seed[1843],seed[2036],seed[3220],seed[3124],seed[1510],seed[1959],seed[2454],seed[859],seed[3474],seed[1550],seed[2179],seed[1143],seed[800],seed[176],seed[2391],seed[1757],seed[3263],seed[1344],seed[647],seed[3398],seed[3379],seed[2231],seed[3213],seed[3527],seed[38],seed[2088],seed[4040],seed[1163],seed[1196],seed[2916],seed[2041],seed[321],seed[31],seed[2676],seed[2548],seed[3438],seed[2025],seed[399],seed[2788],seed[2811],seed[980],seed[1589],seed[2807],seed[465],seed[1853],seed[1902],seed[1019],seed[3488],seed[973],seed[3788],seed[3181],seed[1093],seed[179],seed[679],seed[2137],seed[1248],seed[3400],seed[3901],seed[327],seed[3056],seed[3004],seed[3977],seed[3775],seed[2365],seed[2668],seed[2109],seed[1858],seed[3667],seed[4093],seed[1821],seed[2069],seed[162],seed[2086],seed[2520],seed[493],seed[2337],seed[972],seed[654],seed[1665],seed[545],seed[664],seed[1620],seed[2983],seed[354],seed[595],seed[400],seed[1376],seed[805],seed[1384],seed[3291],seed[1171],seed[2935],seed[1387],seed[1314],seed[3934],seed[4079],seed[1762],seed[1041],seed[310],seed[1036],seed[1198],seed[3482],seed[1353],seed[984],seed[382],seed[223],seed[130],seed[3131],seed[3407],seed[780],seed[1009],seed[2633],seed[1003],seed[1415],seed[876],seed[342],seed[3828],seed[1737],seed[2411],seed[3405],seed[1083],seed[3370],seed[1402],seed[853],seed[1149],seed[2933],seed[2728],seed[444],seed[534],seed[1176],seed[2260],seed[3954],seed[738],seed[1795],seed[1427],seed[2506],seed[983],seed[358],seed[2782],seed[3186],seed[2533],seed[2827],seed[2222],seed[3441],seed[3875],seed[272],seed[3464],seed[1514],seed[1187],seed[3068],seed[3644],seed[2361],seed[978],seed[3548],seed[2999],seed[3745],seed[742],seed[923],seed[2814],seed[2497],seed[3920],seed[70],seed[2977],seed[1808],seed[2080],seed[2071],seed[743],seed[556],seed[3367],seed[2821],seed[4056],seed[2130],seed[1577],seed[2945],seed[1647],seed[626],seed[889],seed[3339],seed[2567],seed[81],seed[1264],seed[340],seed[1379],seed[2403],seed[1385],seed[3969],seed[3294],seed[1796],seed[2981],seed[2015],seed[280],seed[2725],seed[1664],seed[3153],seed[1261],seed[1949],seed[2210],seed[3856],seed[2700],seed[275],seed[3322],seed[955],seed[3242],seed[1408],seed[1776],seed[1400],seed[1260],seed[2435],seed[1989],seed[1416],seed[2398],seed[1390],seed[737],seed[2920],seed[1224],seed[2427],seed[262],seed[1393],seed[15],seed[2597],seed[2372],seed[2318],seed[3361],seed[2483],seed[1883],seed[1106],seed[1477],seed[2924],seed[3661],seed[1226],seed[2755],seed[421],seed[1728],seed[2353],seed[1193],seed[2279],seed[880],seed[412],seed[2525],seed[164],seed[3714],seed[2883],seed[1468],seed[1360],seed[1636],seed[1338],seed[3985],seed[2310],seed[456],seed[1339],seed[3381],seed[1274],seed[3359],seed[2182],seed[2939],seed[2902],seed[767],seed[54],seed[2680],seed[42],seed[602],seed[597],seed[3235],seed[2892],seed[1822],seed[1401],seed[2323],seed[717],seed[2367],seed[831],seed[2049],seed[2993],seed[577],seed[4083],seed[668],seed[3258],seed[625],seed[3401],seed[977],seed[318],seed[3570],seed[1744],seed[1909],seed[908],seed[2370],seed[3557],seed[365],seed[3104],seed[246],seed[462],seed[2949],seed[1317],seed[2666],seed[2004],seed[3063],seed[3026],seed[894],seed[2674],seed[2122],seed[292],seed[1936],seed[2698],seed[4027],seed[1060],seed[3585],seed[1201],seed[1994],seed[1087],seed[2050],seed[1325],seed[424],seed[3731],seed[3274],seed[1194],seed[4088],seed[3463],seed[24],seed[2826],seed[1133],seed[390],seed[2026],seed[2317],seed[3369],seed[1305],seed[2672],seed[2485],seed[2300],seed[2294],seed[2579],seed[985],seed[2505],seed[4045],seed[705],seed[2218],seed[3434],seed[3045],seed[2492],seed[2722],seed[3804],seed[1141],seed[4075],seed[1841],seed[3718],seed[3430],seed[1954],seed[3922],seed[1824],seed[2862],seed[2857],seed[1484],seed[2554],seed[1378],seed[2302],seed[2386],seed[1927],seed[1474],seed[3840],seed[429],seed[3583],seed[159],seed[1673],seed[2248],seed[3574],seed[1667],seed[3368],seed[1835],seed[1061],seed[1210],seed[3457],seed[1492],seed[2641],seed[3330],seed[4016],seed[3481],seed[1605],seed[2019],seed[672],seed[3740],seed[3248],seed[2583],seed[2352],seed[1944],seed[3631],seed[2024],seed[2655],seed[1587],seed[3567],seed[3020],seed[2642],seed[1572],seed[313],seed[1119],seed[4003],seed[830],seed[1945],seed[2268],seed[3619],seed[2032],seed[1575],seed[3394],seed[3766],seed[2192],seed[2211],seed[692],seed[2277],seed[2738],seed[3685],seed[1802],seed[106],seed[2970],seed[3618],seed[2992],seed[2214],seed[1817],seed[3532],seed[2604],seed[4067],seed[2164],seed[1916],seed[2629],seed[3836],seed[953],seed[1663],seed[97],seed[2790],seed[3748],seed[3207],seed[3897],seed[3252],seed[532],seed[3399],seed[1291],seed[3465],seed[932],seed[1350],seed[1644],seed[2127],seed[2224],seed[3284],seed[1321],seed[2747],seed[802],seed[566],seed[916],seed[2275],seed[432],seed[409],seed[1332],seed[1104],seed[1768],seed[1671],seed[3350],seed[2063],seed[2743],seed[2151],seed[904],seed[2720],seed[860],seed[80],seed[1535],seed[700],seed[3891],seed[338],seed[2963],seed[3484],seed[2860],seed[324],seed[1238],seed[813],seed[258],seed[1326],seed[55],seed[1758],seed[2772],seed[600],seed[3756],seed[3929],seed[3940],seed[274],seed[1069],seed[525],seed[2335],seed[3078],seed[473],seed[2091],seed[561],seed[3951],seed[1624],seed[3453],seed[3952],seed[1506],seed[2201],seed[1411],seed[1731],seed[538],seed[603],seed[71],seed[7],seed[2460],seed[2205],seed[3853],seed[1900],seed[2320],seed[773],seed[1188],seed[3133],seed[1983],seed[1423],seed[3173],seed[533],seed[676],seed[4041],seed[2753],seed[245],seed[168],seed[3081],seed[2830],seed[2960],seed[815],seed[2695],seed[1678],seed[2445],seed[3031],seed[520],seed[3072],seed[4064],seed[2582],seed[4037],seed[4055],seed[476],seed[2752],seed[1050],seed[3844],seed[896],seed[2624],seed[1598],seed[1239],seed[3883],seed[2550],seed[482],seed[2379],seed[297],seed[131],seed[2332],seed[2822],seed[2766],seed[641],seed[2219],seed[2756],seed[3955],seed[3102],seed[2566],seed[2220],seed[1372],seed[1056],seed[4046],seed[43],seed[3877],seed[1618],seed[964],seed[3895],seed[2385],seed[3409],seed[2225],seed[3083],seed[1370],seed[1465],seed[3923],seed[2613],seed[2509],seed[2098],seed[3234],seed[2453],seed[1560],seed[1541],seed[2654],seed[1965],seed[433],seed[383],seed[3521],seed[349],seed[463],seed[3306],seed[786],seed[3819],seed[3982],seed[2562],seed[1591],seed[4084],seed[3221],seed[2476],seed[3792],seed[3794],seed[2947],seed[1102],seed[1893],seed[1803],seed[2502],seed[961],seed[920],seed[2298],seed[1156],seed[3467],seed[2486],seed[2750],seed[2552],seed[2420],seed[372],seed[2801],seed[1068],seed[4054],seed[550],seed[631],seed[3495],seed[2481],seed[1232],seed[2659],seed[527],seed[3595],seed[2556],seed[3007],seed[2557],seed[3503],seed[2106],seed[3295],seed[1794],seed[3872],seed[2785],seed[3455],seed[2334],seed[2022],seed[2099],seed[3859],seed[2691],seed[3276],seed[3099],seed[3301],seed[2056],seed[2762],seed[3902],seed[13],seed[3993],seed[1743],seed[3599],seed[593],seed[842],seed[2082],seed[2255],seed[3935],seed[368],seed[1240],seed[753],seed[2479],seed[423],seed[1633],seed[693],seed[552],seed[817],seed[3556],seed[1229],seed[1723],seed[166],seed[2028],seed[1308],seed[2002],seed[1951],seed[790],seed[1948],seed[495],seed[2236],seed[3795],seed[333],seed[1357],seed[1168],seed[3564],seed[2745],seed[3490],seed[2590],seed[2118],seed[2059],seed[3189],seed[136],seed[1209],seed[2072],seed[2459],seed[99],seed[1148],seed[1588],seed[3884],seed[1789],seed[316],seed[388],seed[2794],seed[2033],seed[812],seed[1601],seed[822],seed[1561],seed[852],seed[2784],seed[219],seed[3749],seed[3462],seed[1668],seed[1454],seed[1234],seed[196],seed[3799],seed[732],seed[4011],seed[2396],seed[1355],seed[547],seed[3797],seed[1765],seed[519],seed[2851],seed[3106],seed[1077],seed[2648],seed[2958],seed[2989],seed[3144],seed[3924],seed[3082],seed[1825],seed[1827],seed[384],seed[2769],seed[191],seed[718],seed[2297],seed[962],seed[2416],seed[3577],seed[2816],seed[3832],seed[1760],seed[3148],seed[398],seed[1622],seed[3634],seed[2653],seed[2564],seed[992],seed[1978],seed[1643],seed[1218],seed[1358],seed[841],seed[1581],seed[3609],seed[1130],seed[496],seed[1373],seed[2428],seed[3310],seed[2744],seed[1869],seed[663],seed[3032],seed[1435],seed[2073],seed[3741],seed[3544],seed[1446],seed[640],seed[1862],seed[1786],seed[230],seed[618],seed[2392],seed[3385],seed[3200],seed[588],seed[3192],seed[1710],seed[3265],seed[2046],seed[2390],seed[677],seed[3108],seed[1798],seed[1154],seed[857],seed[847],seed[367],seed[330],seed[374],seed[3890],seed[210],seed[2940],seed[2684],seed[3991],seed[1329],seed[1159],seed[3814],seed[891],seed[1943],seed[2805],seed[1775],seed[3972],seed[3043],seed[1684],seed[406],seed[3348],seed[517],seed[312],seed[3687],seed[3468],seed[2560],seed[3960],seed[466],seed[3046],seed[574],seed[3755],seed[791],seed[1582],seed[3860],seed[2682],seed[1553],seed[2336],seed[1137],seed[1230],seed[2842],seed[2121],seed[617],seed[804],seed[2200],seed[1650],seed[715],seed[2657],seed[3497],seed[2893],seed[3296],seed[2596],seed[531],seed[2809],seed[143],seed[3170],seed[1928],seed[1654],seed[2124],seed[4070],seed[3927],seed[3805],seed[2957],seed[322],seed[1430],seed[356],seed[397],seed[119],seed[3600],seed[1000],seed[3944],seed[252],seed[1666],seed[788],seed[2434],seed[3431],seed[1896],seed[1086],seed[1250],seed[3387],seed[1791],seed[1303],seed[3781],seed[1584],seed[2344],seed[2953],seed[1412],seed[3601],seed[1819],seed[2946],seed[497],seed[3445],seed[1691],seed[1558],seed[2995],seed[3347],seed[607],seed[3966],seed[1689],seed[951],seed[558],seed[3143],seed[487],seed[4058],seed[1070],seed[2507],seed[2727],seed[154],seed[1351],seed[3916],seed[2938],seed[1312],seed[2395],seed[1999],seed[1183],seed[170],seed[56],seed[460],seed[75],seed[2456],seed[2311],seed[2010],seed[914],seed[10],seed[3997],seed[688],seed[845],seed[3000],seed[4013],seed[3695],seed[2215],seed[2290],seed[2994],seed[3341],seed[843],seed[1868],seed[3911],seed[3053],seed[709],seed[121],seed[2976],seed[3215],seed[295],seed[2239],seed[1085],seed[1029],seed[2898],seed[2662],seed[227],seed[645],seed[2894],seed[1679],seed[77],seed[1206],seed[1147],seed[591],seed[3270],seed[2911],seed[3416],seed[1276],seed[350],seed[2491],seed[2915],seed[739],seed[2884],seed[1814],seed[2014],seed[2937],seed[255],seed[1464],seed[3713],seed[2796],seed[2308],seed[2227],seed[385],seed[4035],seed[1310],seed[781],seed[1144],seed[1769],seed[2415],seed[567],seed[4094],seed[1640],seed[1960],seed[68],seed[2440],seed[1213],seed[187],seed[326],seed[869],seed[2917],seed[2394],seed[3404],seed[1409],seed[884],seed[2645],seed[502],seed[2797],seed[3870],seed[257],seed[3703],seed[3206],seed[2038],seed[1440],seed[452],seed[2735],seed[3679],seed[1242],seed[3514],seed[1192],seed[3803],seed[3621],seed[704],seed[1501],seed[1603],seed[562],seed[3889],seed[171],seed[1991],seed[3500],seed[2663],seed[3605],seed[3277],seed[2433],seed[234],seed[3617],seed[766],seed[4029],seed[2694],seed[298],seed[2155],seed[1146],seed[1534],seed[1391],seed[427],seed[3727],seed[596],seed[1225],seed[2226],seed[2897],seed[3364],seed[1755],seed[3635],seed[1472],seed[3719],seed[3636],seed[756],seed[2321],seed[1251],seed[2383],seed[3217],seed[1958],seed[1398],seed[2715],seed[1420],seed[3677],seed[2177],seed[1217],seed[1611],seed[3425],seed[3435],seed[416],seed[2586],seed[3700],seed[3938],seed[3823],seed[1457],seed[3149],seed[1328],seed[2358],seed[1257],seed[1051],seed[3150],seed[1565],seed[3062],seed[3470],seed[1109],seed[1418],seed[2402],seed[2854],seed[3121],seed[1216],seed[1736],seed[3334],seed[2055],seed[1612],seed[1854],seed[4006],seed[1],seed[3864],seed[2262],seed[3758],seed[864],seed[819],seed[3898],seed[1641],seed[4044],seed[2825],seed[2257],seed[2053],seed[2085],seed[2577],seed[1121],seed[1190],seed[1236],seed[1992],seed[320],seed[353],seed[2671],seed[635],seed[2223],seed[2430],seed[644],seed[3298],seed[3672],seed[3204],seed[3907],seed[152],seed[3038],seed[3673],seed[1030],seed[3613],seed[956],seed[1521],seed[2882],seed[3224],seed[3646],seed[2076],seed[2644],seed[2304],seed[165],seed[2996],seed[485],seed[3432],seed[1837],seed[1311],seed[2446],seed[724],seed[513],seed[1963],seed[3774],seed[2347],seed[3100],seed[1269],seed[1811],seed[3163],seed[3125],seed[2207],seed[180],seed[3682],seed[377],seed[1480],seed[105],seed[2833],seed[1460],seed[3946],seed[3127],seed[1204],seed[2504],seed[2852],seed[3690],seed[3380],seed[20],seed[3833],seed[3534],seed[1523],seed[3625],seed[5],seed[1164],seed[939],seed[1635],seed[2757],seed[3592],seed[2061],seed[1766],seed[1333],seed[3262],seed[2763],seed[1773],seed[3624],seed[3620],seed[2609],seed[1846],seed[2656],seed[638],seed[3563],seed[35],seed[3251],seed[730],seed[2443],seed[468],seed[634],seed[335],seed[3185],seed[315],seed[2532],seed[3172],seed[8],seed[3581],seed[2461],seed[3671],seed[2016],seed[145],seed[1745],seed[1132],seed[483],seed[606],seed[621],seed[1369],seed[464],seed[1695],seed[2518],seed[3632],seed[3704],seed[331],seed[835],seed[3442],seed[690],seed[765],seed[156],seed[391],seed[1838],seed[2956],seed[1848],seed[3806],seed[1533],seed[1675],seed[3588],seed[2716],seed[243],seed[2626],seed[49],seed[2867],seed[3243],seed[643],seed[3487],seed[686],seed[3706],seed[604],seed[2547],seed[3344],seed[402],seed[2943],seed[528],seed[3414],seed[4033],seed[2627],seed[253],seed[3863],seed[993],seed[3309],seed[1968],seed[134],seed[2985],seed[1284],seed[3539],seed[1175],seed[3021],seed[211],seed[1683],seed[355],seed[453],seed[4032],seed[1122],seed[794],seed[446],seed[3249],seed[2423],seed[699],seed[378],seed[3917],seed[3879],seed[810],seed[2664],seed[1017],seed[1870],seed[3835],seed[1716],seed[3443],seed[2647],seed[1545],seed[670],seed[1424],seed[2699],seed[129],seed[1599],seed[2147],seed[3132],seed[4026],seed[1607],seed[2194],seed[3678],seed[3461],seed[1431],seed[2351],seed[2864],seed[1428],seed[684],seed[1895],seed[2871],seed[3639],seed[3862],seed[478],seed[2831],seed[2208],seed[2887],seed[2693],seed[770],seed[899],seed[2839],seed[46],seed[2503],seed[1380],seed[2665],seed[1966],seed[1422],seed[2040],seed[1897],seed[2345],seed[2623],seed[3029],seed[1235],seed[2880],seed[197],seed[3420],seed[2510],seed[1924],seed[1266],seed[1025],seed[1842],seed[3992],seed[712],seed[2602],seed[2606],seed[1865],seed[2203],seed[892],seed[504],seed[1705],seed[877],seed[3228],seed[64],seed[2966],seed[3522],seed[2449],seed[2499],seed[573],seed[1935],seed[2603],seed[3202],seed[306],seed[461],seed[431],seed[722],seed[2705],seed[3820],seed[3928],seed[1890],seed[2612],seed[3787],seed[963],seed[3332],seed[3233],seed[1833],seed[2760],seed[1478],seed[1878],seed[3329],seed[1756],seed[2013],seed[214],seed[265],seed[975],seed[1139],seed[3103],seed[1455],seed[582],seed[807],seed[2789],seed[389],seed[3239],seed[3061],seed[4],seed[1300],seed[2330],seed[2424],seed[3041],seed[3337],seed[710],seed[2009],seed[777],seed[1810],seed[3752],seed[2465],seed[2931],seed[3049],seed[3071],seed[414],seed[2045],seed[2929],seed[785],seed[3650],seed[675],seed[2284],seed[101],seed[707],seed[1103],seed[2114],seed[3093],seed[1334],seed[3473],seed[23],seed[3184],seed[1397],seed[3389],seed[1672],seed[3926],seed[2142],seed[3722],seed[3036],seed[2584],seed[422],seed[3878],seed[205],seed[2413],seed[3384],seed[1770],seed[3770],seed[968],seed[3717],seed[249],seed[2859],seed[314],seed[1522],seed[2683],seed[529],seed[3151],seed[2261],seed[3665],seed[936],seed[854],seed[4025],seed[4051],seed[172],seed[1826],seed[1114],seed[970],seed[2517],seed[3074],seed[1638],seed[1986],seed[299],seed[3763],seed[1487],seed[1911],seed[2338],seed[4062],seed[3762],seed[1552],seed[273],seed[225],seed[1436],seed[938],seed[2442],seed[3223],seed[913],seed[2293],seed[2247],seed[2542],seed[999],seed[3304],seed[945],seed[3518],seed[1105],seed[2163],seed[2622],seed[1659],seed[3012],seed[598],seed[58],seed[2314],seed[636],seed[1805],seed[3655],seed[2614],seed[123],seed[3777],seed[541],seed[967],seed[4060]}),
        .cross_prob(cross_prob),
        .codeword(codeword13),
        .received(received13)
        );
    
    bsc bsc14(
        .clk(clk),
        .reset(reset),
        .seed({seed[2718],seed[1655],seed[1349],seed[2651],seed[2271],seed[1920],seed[2133],seed[3033],seed[1147],seed[3493],seed[3143],seed[3813],seed[1282],seed[965],seed[2138],seed[3855],seed[1779],seed[2163],seed[3446],seed[1444],seed[109],seed[1414],seed[2943],seed[2341],seed[1598],seed[2033],seed[628],seed[2861],seed[1758],seed[3119],seed[2265],seed[2479],seed[3910],seed[271],seed[1139],seed[1006],seed[2361],seed[1930],seed[979],seed[91],seed[1843],seed[3617],seed[3190],seed[993],seed[2217],seed[2001],seed[3822],seed[873],seed[1510],seed[1924],seed[522],seed[612],seed[777],seed[1891],seed[757],seed[2219],seed[3352],seed[1218],seed[1348],seed[3199],seed[3260],seed[1576],seed[2537],seed[3373],seed[2956],seed[3018],seed[1462],seed[2522],seed[1820],seed[3148],seed[3688],seed[647],seed[3264],seed[2481],seed[1481],seed[365],seed[1938],seed[1752],seed[1411],seed[2004],seed[65],seed[2470],seed[4090],seed[3276],seed[501],seed[312],seed[3236],seed[939],seed[1571],seed[3080],seed[1525],seed[926],seed[3285],seed[1984],seed[764],seed[3680],seed[1328],seed[1251],seed[2516],seed[2258],seed[3667],seed[879],seed[872],seed[3379],seed[2659],seed[3126],seed[1508],seed[3381],seed[90],seed[1677],seed[2693],seed[3777],seed[7],seed[3610],seed[1181],seed[3637],seed[3189],seed[2740],seed[1352],seed[1237],seed[1198],seed[2419],seed[606],seed[14],seed[94],seed[1682],seed[2630],seed[2365],seed[1704],seed[2488],seed[1177],seed[2600],seed[2679],seed[1059],seed[914],seed[1472],seed[3521],seed[1199],seed[3991],seed[1337],seed[1153],seed[2552],seed[2994],seed[1267],seed[4016],seed[281],seed[3696],seed[2746],seed[421],seed[2327],seed[3536],seed[1997],seed[12],seed[3640],seed[2181],seed[3170],seed[294],seed[665],seed[1724],seed[517],seed[2476],seed[2967],seed[2503],seed[568],seed[1273],seed[2698],seed[3862],seed[3556],seed[2624],seed[1882],seed[1841],seed[592],seed[3642],seed[3205],seed[2287],seed[3280],seed[2373],seed[1538],seed[3097],seed[4051],seed[2836],seed[2834],seed[431],seed[2399],seed[3339],seed[2773],seed[1769],seed[2420],seed[3716],seed[1357],seed[2526],seed[3413],seed[1255],seed[384],seed[637],seed[713],seed[1464],seed[27],seed[3408],seed[135],seed[3055],seed[3215],seed[537],seed[2964],seed[3830],seed[2034],seed[383],seed[2066],seed[3449],seed[3477],seed[3098],seed[3090],seed[1520],seed[3155],seed[1903],seed[3824],seed[1913],seed[805],seed[1660],seed[656],seed[161],seed[3990],seed[661],seed[3041],seed[3917],seed[2543],seed[728],seed[1026],seed[2121],seed[1130],seed[3618],seed[3258],seed[2549],seed[268],seed[1917],seed[2412],seed[1263],seed[8],seed[802],seed[307],seed[2762],seed[1766],seed[3208],seed[2132],seed[3913],seed[1887],seed[3237],seed[1597],seed[604],seed[2865],seed[3432],seed[1961],seed[3766],seed[1505],seed[3218],seed[166],seed[120],seed[3300],seed[3374],seed[574],seed[538],seed[2665],seed[1032],seed[460],seed[3178],seed[2179],seed[2395],seed[1308],seed[652],seed[591],seed[2973],seed[617],seed[3593],seed[1848],seed[744],seed[3038],seed[3393],seed[704],seed[2821],seed[1854],seed[1523],seed[1201],seed[751],seed[1384],seed[2177],seed[3972],seed[2366],seed[1304],seed[1565],seed[3054],seed[2246],seed[413],seed[3816],seed[3590],seed[4026],seed[689],seed[2619],seed[1389],seed[500],seed[3282],seed[3130],seed[1594],seed[437],seed[916],seed[3011],seed[3865],seed[2403],seed[3516],seed[2962],seed[1974],seed[1128],seed[3158],seed[1784],seed[105],seed[1729],seed[3962],seed[1764],seed[3454],seed[2997],seed[1089],seed[1129],seed[718],seed[2433],seed[2013],seed[1585],seed[1686],seed[3946],seed[2256],seed[3444],seed[745],seed[2417],seed[29],seed[1725],seed[1787],seed[3140],seed[1007],seed[2368],seed[1477],seed[1539],seed[1794],seed[2996],seed[148],seed[3501],seed[2839],seed[3100],seed[2780],seed[1928],seed[3875],seed[2255],seed[2761],seed[2371],seed[302],seed[3682],seed[2618],seed[638],seed[1950],seed[723],seed[3572],seed[104],seed[4052],seed[1034],seed[385],seed[1061],seed[2335],seed[3240],seed[2176],seed[3228],seed[1722],seed[2095],seed[4003],seed[2782],seed[531],seed[1042],seed[3058],seed[3641],seed[2697],seed[2979],seed[382],seed[904],seed[84],seed[4070],seed[3294],seed[4009],seed[1781],seed[219],seed[3936],seed[2505],seed[2827],seed[284],seed[2666],seed[4005],seed[953],seed[3878],seed[2980],seed[1625],seed[3136],seed[1424],seed[511],seed[934],seed[3817],seed[3230],seed[1790],seed[836],seed[414],seed[1159],seed[3753],seed[3835],seed[3284],seed[1833],seed[2615],seed[3006],seed[3540],seed[1618],seed[3635],seed[3082],seed[3067],seed[1207],seed[1761],seed[3845],seed[1912],seed[1735],seed[3971],seed[1964],seed[1829],seed[3951],seed[1203],seed[3425],seed[110],seed[3307],seed[2143],seed[1617],seed[75],seed[2289],seed[3989],seed[3928],seed[2941],seed[454],seed[2506],seed[2447],seed[3330],seed[3639],seed[2146],seed[278],seed[308],seed[567],seed[554],seed[2750],seed[1688],seed[2885],seed[2038],seed[4014],seed[2749],seed[2947],seed[1856],seed[2915],seed[703],seed[1527],seed[3278],seed[2092],seed[1972],seed[3698],seed[3324],seed[1710],seed[2079],seed[425],seed[440],seed[206],seed[2111],seed[707],seed[4031],seed[2422],seed[1246],seed[3040],seed[3418],seed[1355],seed[3767],seed[851],seed[3726],seed[1036],seed[3973],seed[2064],seed[1316],seed[2999],seed[2873],seed[1786],seed[2633],seed[3654],seed[2021],seed[748],seed[597],seed[3009],seed[1692],seed[131],seed[3206],seed[2431],seed[1706],seed[2931],seed[528],seed[2350],seed[3792],seed[932],seed[1120],seed[1734],seed[898],seed[3160],seed[357],seed[2654],seed[903],seed[2290],seed[3281],seed[3725],seed[1543],seed[3029],seed[253],seed[3077],seed[1663],seed[2667],seed[2877],seed[215],seed[2923],seed[633],seed[3941],seed[2444],seed[927],seed[806],seed[1166],seed[1838],seed[601],seed[2691],seed[890],seed[2660],seed[2108],seed[2547],seed[2270],seed[3226],seed[1367],seed[185],seed[3219],seed[125],seed[60],seed[3386],seed[2778],seed[1522],seed[3524],seed[2957],seed[2316],seed[2074],seed[783],seed[840],seed[3378],seed[2484],seed[130],seed[1405],seed[2220],seed[1956],seed[349],seed[3626],seed[2497],seed[3305],seed[2105],seed[1172],seed[2715],seed[2527],seed[350],seed[2156],seed[328],seed[2449],seed[1380],seed[1802],seed[2360],seed[4019],seed[471],seed[406],seed[2813],seed[797],seed[2596],seed[158],seed[122],seed[3351],seed[1588],seed[1014],seed[180],seed[493],seed[1979],seed[3474],seed[4048],seed[313],seed[3153],seed[721],seed[3820],seed[2154],seed[96],seed[2791],seed[1043],seed[4006],seed[2427],seed[2211],seed[3052],seed[1814],seed[167],seed[1926],seed[648],seed[3580],seed[3288],seed[3037],seed[237],seed[3229],seed[2981],seed[3472],seed[2134],seed[2717],seed[121],seed[2195],seed[2560],seed[321],seed[3814],seed[182],seed[2758],seed[3883],seed[509],seed[2644],seed[2607],seed[2169],seed[3560],seed[1876],seed[20],seed[404],seed[828],seed[945],seed[174],seed[2508],seed[147],seed[825],seed[2533],seed[2261],seed[1792],seed[2765],seed[3597],seed[544],seed[1503],seed[1236],seed[2755],seed[543],seed[3712],seed[99],seed[3473],seed[1487],seed[3988],seed[1134],seed[2763],seed[1416],seed[3577],seed[4000],seed[1229],seed[552],seed[3721],seed[1743],seed[3089],seed[2187],seed[1087],seed[1124],seed[2523],seed[2472],seed[2022],seed[286],seed[98],seed[4035],seed[1874],seed[1708],seed[463],seed[2230],seed[176],seed[1002],seed[3411],seed[919],seed[2656],seed[822],seed[583],seed[782],seed[2393],seed[1277],seed[790],seed[1265],seed[3396],seed[2262],seed[881],seed[2223],seed[3749],seed[3841],seed[1826],seed[3387],seed[3921],seed[4037],seed[2385],seed[2392],seed[3670],seed[632],seed[3863],seed[513],seed[1537],seed[3484],seed[2482],seed[2952],seed[3558],seed[395],seed[1817],seed[1458],seed[423],seed[1433],seed[2315],seed[870],seed[126],seed[1687],seed[2298],seed[2905],seed[5],seed[1716],seed[2291],seed[3608],seed[3275],seed[1528],seed[2390],seed[3860],seed[265],seed[1593],seed[1944],seed[0],seed[2858],seed[1546],seed[288],seed[2308],seed[1100],seed[181],seed[1855],seed[3856],seed[1497],seed[2218],seed[3809],seed[3162],seed[2535],seed[2018],seed[1209],seed[2669],seed[407],seed[2539],seed[3684],seed[3853],seed[2306],seed[157],seed[1023],seed[1774],seed[1737],seed[3554],seed[856],seed[2463],seed[1090],seed[716],seed[2672],seed[1985],seed[1257],seed[3195],seed[3507],seed[3061],seed[3899],seed[2436],seed[1581],seed[3919],seed[2362],seed[3397],seed[2090],seed[2297],seed[3960],seed[1064],seed[1278],seed[2907],seed[2948],seed[3429],seed[3065],seed[3615],seed[2023],seed[2515],seed[3581],seed[2151],seed[175],seed[2448],seed[2793],seed[3812],seed[410],seed[2029],seed[3401],seed[3837],seed[762],seed[3606],seed[2716],seed[4057],seed[1286],seed[2052],seed[959],seed[3966],seed[603],seed[2728],seed[3548],seed[848],seed[865],seed[1048],seed[621],seed[277],seed[3768],seed[2859],seed[3594],seed[2234],seed[459],seed[2369],seed[2601],seed[3481],seed[3075],seed[640],seed[759],seed[332],seed[4013],seed[3673],seed[690],seed[4010],seed[3685],seed[82],seed[149],seed[1154],seed[1919],seed[2880],seed[3326],seed[267],seed[2807],seed[2326],seed[1501],seed[1805],seed[3629],seed[774],seed[4032],seed[521],seed[1270],seed[2511],seed[4073],seed[2178],seed[272],seed[818],seed[3166],seed[1951],seed[1310],seed[4007],seed[3665],seed[3415],seed[3889],seed[3131],seed[4002],seed[247],seed[2490],seed[3675],seed[455],seed[838],seed[3069],seed[949],seed[2838],seed[2707],seed[1183],seed[364],seed[3949],seed[2845],seed[3539],seed[3464],seed[2816],seed[3471],seed[1850],seed[2115],seed[264],seed[2574],seed[1696],seed[3181],seed[3430],seed[129],seed[4047],seed[3791],seed[666],seed[2123],seed[244],seed[3801],seed[670],seed[920],seed[1858],seed[1999],seed[1504],seed[1359],seed[1379],seed[2814],seed[2922],seed[1863],seed[2673],seed[3914],seed[266],seed[2280],seed[2235],seed[3360],seed[3727],seed[2440],seed[3839],seed[3492],seed[389],seed[1131],seed[2823],seed[518],seed[2453],seed[4075],seed[3745],seed[2008],seed[758],seed[2507],seed[361],seed[1605],seed[1676],seed[896],seed[588],seed[112],seed[2128],seed[2810],seed[2846],seed[3690],seed[34],seed[1822],seed[1506],seed[1670],seed[3840],seed[1055],seed[3161],seed[143],seed[3355],seed[1008],seed[3515],seed[1816],seed[3699],seed[33],seed[3347],seed[3505],seed[171],seed[231],seed[859],seed[2592],seed[1895],seed[2971],seed[3269],seed[2863],seed[3296],seed[1419],seed[769],seed[1213],seed[1327],seed[2227],seed[4017],seed[3409],seed[1610],seed[3895],seed[1775],seed[846],seed[2048],seed[3013],seed[2245],seed[676],seed[664],seed[2175],seed[2257],seed[3705],seed[2955],seed[3405],seed[426],seed[1275],seed[3969],seed[2379],seed[1215],seed[709],seed[381],seed[1493],seed[1910],seed[651],seed[2870],seed[275],seed[3701],seed[1170],seed[2414],seed[2556],seed[453],seed[3672],seed[529],seed[964],seed[204],seed[2058],seed[2895],seed[3894],seed[352],seed[1496],seed[2323],seed[2803],seed[784],seed[1550],seed[3297],seed[114],seed[826],seed[639],seed[921],seed[69],seed[1434],seed[1473],seed[3335],seed[3873],seed[1762],seed[2231],seed[1853],seed[2978],seed[1544],seed[2963],seed[3785],seed[2078],seed[1322],seed[3761],seed[297],seed[2321],seed[733],seed[958],seed[4067],seed[771],seed[2221],seed[1827],seed[2239],seed[2016],seed[3354],seed[3589],seed[1712],seed[3116],seed[1992],seed[2404],seed[2467],seed[1070],seed[3030],seed[3486],seed[1443],seed[658],seed[1630],seed[3514],seed[1902],seed[3293],seed[735],seed[358],seed[2478],seed[2712],seed[134],seed[2454],seed[594],seed[616],seed[823],seed[3453],seed[2721],seed[1076],seed[240],seed[3087],seed[245],seed[3943],seed[2370],seed[1842],seed[1394],seed[235],seed[1016],seed[2835],seed[1499],seed[839],seed[1371],seed[1083],seed[2713],seed[1217],seed[3213],seed[52],seed[3020],seed[2595],seed[292],seed[2710],seed[1921],seed[3341],seed[2338],seed[3487],seed[1939],seed[1418],seed[2983],seed[1723],seed[3634],seed[2599],seed[2376],seed[907],seed[3068],seed[2450],seed[1],seed[2992],seed[1693],seed[971],seed[2046],seed[3081],seed[1574],seed[1960],seed[572],seed[2510],seed[1234],seed[2700],seed[3246],seed[2501],seed[996],seed[1620],seed[3833],seed[795],seed[2685],seed[2277],seed[1513],seed[331],seed[2893],seed[3553],seed[1552],seed[1085],seed[3321],seed[3694],seed[3920],seed[480],seed[1179],seed[3198],seed[2896],seed[1141],seed[1634],seed[1763],seed[3295],seed[3623],seed[3248],seed[1216],seed[3057],seed[3245],seed[3366],seed[3123],seed[1661],seed[1260],seed[2041],seed[1088],seed[3599],seed[1629],seed[1377],seed[3436],seed[843],seed[2653],seed[813],seed[577],seed[283],seed[1832],seed[1953],seed[1241],seed[3191],seed[3380],seed[169],seed[3107],seed[2632],seed[320],seed[319],seed[1212],seed[2465],seed[448],seed[3834],seed[386],seed[355],seed[2076],seed[1649],seed[187],seed[3600],seed[615],seed[3700],seed[1163],seed[809],seed[2932],seed[1290],seed[863],seed[1884],seed[3573],seed[3438],seed[2590],seed[2437],seed[3825],seed[2611],seed[433],seed[645],seed[2011],seed[1906],seed[3182],seed[992],seed[2789],seed[598],seed[3095],seed[2631],seed[3252],seed[546],seed[2408],seed[3103],seed[2689],seed[2593],seed[2864],seed[623],seed[374],seed[3740],seed[2645],seed[1969],seed[3194],seed[1797],seed[1904],seed[3337],seed[3986],seed[3729],seed[47],seed[1640],seed[683],seed[3645],seed[1783],seed[3124],seed[1400],seed[3406],seed[197],seed[3203],seed[860],seed[833],seed[1295],seed[1536],seed[3186],seed[3806],seed[1828],seed[2616],seed[669],seed[2891],seed[3154],seed[3202],seed[470],seed[956],seed[89],seed[2899],seed[2609],seed[2324],seed[2826],seed[2387],seed[2898],seed[291],seed[941],seed[3746],seed[1456],seed[2317],seed[378],seed[2843],seed[444],seed[3327],seed[2206],seed[3995],seed[3728],seed[3403],seed[504],seed[3660],seed[620],seed[1314],seed[1778],seed[2777],seed[4015],seed[80],seed[2039],seed[1350],seed[3596],seed[724],seed[634],seed[2486],seed[41],seed[1081],seed[2459],seed[3965],seed[2068],seed[1857],seed[2005],seed[2065],seed[2259],seed[1809],seed[1202],seed[2538],seed[446],seed[1045],seed[429],seed[1249],seed[2544],seed[557],seed[2725],seed[902],seed[611],seed[1301],seed[2568],seed[2736],seed[1987],seed[832],seed[394],seed[1342],seed[3249],seed[2037],seed[1364],seed[2944],seed[2796],seed[224],seed[1027],seed[553],seed[2563],seed[1633],seed[3157],seed[3592],seed[1345],seed[2180],seed[1937],seed[2456],seed[2714],seed[2435],seed[2352],seed[3538],seed[533],seed[2771],seed[322],seed[2167],seed[1066],seed[438],seed[3882],seed[3537],seed[2995],seed[1541],seed[227],seed[2288],seed[3268],seed[827],seed[3666],seed[1005],seed[1341],seed[1127],seed[3723],seed[299],seed[753],seed[702],seed[2402],seed[1022],seed[1266],seed[481],seed[899],seed[3021],seed[2901],seed[1907],seed[259],seed[1340],seed[1180],seed[2060],seed[1830],seed[2168],seed[329],seed[1720],seed[68],seed[2702],seed[1185],seed[1835],seed[3361],seed[464],seed[3783],seed[3110],seed[3849],seed[3368],seed[37],seed[3513],seed[581],seed[749],seed[2149],seed[2910],seed[3846],seed[3784],seed[2102],seed[2426],seed[3927],seed[1467],seed[1475],seed[3437],seed[432],seed[401],seed[2764],seed[368],seed[309],seed[3836],seed[3713],seed[1654],seed[59],seed[97],seed[3083],seed[1892],seed[2745],seed[1518],seed[3650],seed[2131],seed[457],seed[2682],seed[3025],seed[3479],seed[1671],seed[2489],seed[77],seed[2112],seed[2344],seed[711],seed[2760],seed[1507],seed[1911],seed[3359],seed[3102],seed[2043],seed[3747],seed[391],seed[3942],seed[3072],seed[1426],seed[1235],seed[697],seed[1806],seed[2358],seed[3490],seed[915],seed[258],seed[1200],seed[2868],seed[1148],seed[1437],seed[1511],seed[514],seed[2455],seed[417],seed[877],seed[1041],seed[177],seed[2583],seed[788],seed[1227],seed[3674],seed[1665],seed[1867],seed[2844],seed[2951],seed[3775],seed[1190],seed[1698],seed[2965],seed[127],seed[1001],seed[3510],seed[3008],seed[3715],seed[2770],seed[4065],seed[145],seed[1936],seed[869],seed[151],seed[3903],seed[1749],seed[1846],seed[2798],seed[492],seed[2430],seed[844],seed[495],seed[800],seed[910],seed[3506],seed[1674],seed[2812],seed[3096],seed[969],seed[2743],seed[3050],seed[857],seed[1033],seed[663],seed[3693],seed[3063],seed[155],seed[2164],seed[1169],seed[1356],seed[3261],seed[1450],seed[3497],seed[2418],seed[2850],seed[50],seed[2117],seed[4039],seed[3758],seed[1877],seed[1715],seed[324],seed[972],seed[1645],seed[1178],seed[373],seed[1488],seed[3048],seed[2055],seed[1427],seed[26],seed[379],seed[808],seed[1440],seed[4084],seed[2421],seed[1140],seed[2976],seed[3823],seed[2559],seed[3522],seed[2640],seed[1868],seed[2818],seed[3016],seed[3176],seed[1900],seed[478],seed[654],seed[1370],seed[1714],seed[3821],seed[1412],seed[3980],seed[3452],seed[2988],seed[1113],seed[3710],seed[786],seed[649],seed[3333],seed[4080],seed[883],seed[2283],seed[1932],seed[3854],seed[1922],seed[3706],seed[3212],seed[3099],seed[1143],seed[3085],seed[629],seed[842],seed[3101],seed[3868],seed[1927],seed[961],seed[2364],seed[2495],seed[3983],seed[86],seed[3256],seed[2423],seed[3638],seed[4041],seed[1390],seed[252],seed[1871],seed[1259],seed[1847],seed[4030],seed[1648],seed[342],seed[2542],seed[655],seed[878],seed[2786],seed[3384],seed[3552],seed[3891],seed[1431],seed[2212],seed[1455],seed[1878],seed[300],seed[2639],seed[2614],seed[3350],seed[3168],seed[2116],seed[2572],seed[1554],seed[1108],seed[3483],seed[3221],seed[203],seed[1478],seed[92],seed[950],seed[1553],seed[3851],seed[1062],seed[387],seed[787],seed[1012],seed[1726],seed[2329],seed[3736],seed[1274],seed[3496],seed[3367],seed[726],seed[3717],seed[3754],seed[1053],seed[3652],seed[1616],seed[424],seed[3211],seed[419],seed[2792],seed[1524],seed[3024],seed[503],seed[3431],seed[276],seed[1192],seed[2851],seed[2819],seed[2558],seed[3542],seed[3533],seed[3201],seed[137],seed[2494],seed[1373],seed[2741],seed[36],seed[3056],seed[2986],seed[2309],seed[399],seed[390],seed[867],seed[3764],seed[2555],seed[3108],seed[213],seed[2357],seed[2445],seed[2902],seed[2781],seed[2363],seed[3074],seed[2340],seed[761],seed[2513],seed[2040],seed[1718],seed[3789],seed[229],seed[1395],seed[2929],seed[2575],seed[3343],seed[2954],seed[1941],seed[855],seed[3826],seed[3940],seed[678],seed[2442],seed[3465],seed[3036],seed[3689],seed[2610],seed[696],seed[3730],seed[3287],seed[436],seed[2017],seed[2030],seed[549],seed[816],seed[2657],seed[3861],seed[1568],seed[1562],seed[434],seed[2135],seed[1592],seed[2401],seed[251],seed[2356],seed[1705],seed[376],seed[306],seed[2215],seed[2726],seed[2477],seed[3028],seed[3714],seed[1287],seed[1311],seed[3267],seed[274],seed[1430],seed[226],seed[2010],seed[502],seed[1482],seed[991],seed[2160],seed[610],seed[3504],seed[2293],seed[3997],seed[260],seed[1759],seed[3755],seed[3489],seed[1560],seed[3263],seed[173],seed[2140],seed[1285],seed[2587],seed[801],seed[2471],seed[1545],seed[2950],seed[273],seed[635],seed[35],seed[3111],seed[363],seed[2388],seed[3531],seed[3773],seed[2110],seed[241],seed[3117],seed[1897],seed[2779],seed[427],seed[3400],seed[687],seed[1767],seed[1193],seed[569],seed[2382],seed[2330],seed[794],seed[3372],seed[785],seed[1746],seed[681],seed[3984],seed[3896],seed[3901],seed[3994],seed[1567],seed[1044],seed[3079],seed[325],seed[2534],seed[1619],seed[1711],seed[1879],seed[326],seed[2553],seed[1232],seed[1751],seed[2748],seed[952],seed[483],seed[819],seed[507],seed[2057],seed[79],seed[2020],seed[1451],seed[1777],seed[2093],seed[1245],seed[1849],seed[776],seed[3898],seed[2084],seed[3273],seed[876],seed[738],seed[1191],seed[354],seed[1901],seed[2451],seed[804],seed[3325],seed[1396],seed[76],seed[3549],seed[3187],seed[2487],seed[1840],seed[3047],seed[2620],seed[1942],seed[4078],seed[3532],seed[1547],seed[4024],seed[614],seed[922],seed[2801],seed[3105],seed[2564],seed[2841],seed[3338],seed[3760],seed[2424],seed[817],seed[1258],seed[1078],seed[3466],seed[3576],seed[1461],seed[1300],seed[186],seed[1925],seed[3907],seed[3462],seed[163],seed[2808],seed[330],seed[798],seed[3291],seed[803],seed[3708],seed[3336],seed[2696],seed[1402],seed[3525],seed[3979],seed[3671],seed[3850],seed[183],seed[1933],seed[1952],seed[2541],seed[2342],seed[2622],seed[2594],seed[3259],seed[695],seed[1335],seed[2213],seed[2145],seed[2848],seed[1521],seed[3864],seed[3423],seed[1292],seed[2322],seed[1152],seed[2753],seed[1470],seed[987],seed[3751],seed[411],seed[1065],seed[345],seed[1793],seed[1291],seed[1293],seed[2222],seed[2884],seed[2975],seed[2443],seed[3383],seed[2768],seed[2049],seed[3053],seed[1247],seed[1404],seed[3551],seed[590],seed[831],seed[506],seed[409],seed[1406],seed[3495],seed[3686],seed[555],seed[1358],seed[4082],seed[1220],seed[1151],seed[344],seed[2158],seed[78],seed[1142],seed[4068],seed[2514],seed[2263],seed[754],seed[375],seed[3209],seed[1063],seed[1176],seed[1584],seed[1423],seed[449],seed[3315],seed[208],seed[2059],seed[3842],seed[1347],seed[3316],seed[3439],seed[2069],seed[2822],seed[3470],seed[102],seed[249],seed[541],seed[3426],seed[3961],seed[1319],seed[3445],seed[2304],seed[1570],seed[3344],seed[3559],seed[2272],seed[2407],seed[1360],seed[1004],seed[2678],seed[262],seed[1731],seed[3948],seed[1614],seed[2927],seed[3142],seed[1020],seed[2464],seed[1339],seed[2968],seed[3857],seed[1174],seed[4056],seed[4036],seed[2268],seed[136],seed[1155],seed[3370],seed[742],seed[2674],seed[3322],seed[743],seed[712],seed[4061],seed[2809],seed[1559],seed[1557],seed[3217],seed[2044],seed[3032],seed[1336],seed[362],seed[3697],seed[1975],seed[1949],seed[2229],seed[2378],seed[2075],seed[980],seed[3779],seed[3014],seed[2007],seed[3695],seed[3603],seed[3923],seed[2663],seed[1317],seed[3459],seed[1946],seed[3547],seed[3109],seed[195],seed[3238],seed[2284],seed[1401],seed[2498],seed[1851],seed[3262],seed[2091],seed[2087],seed[3681],seed[731],seed[10],seed[201],seed[1608],seed[1866],seed[2739],seed[2990],seed[2279],seed[2249],seed[3739],seed[2207],seed[1821],seed[3141],seed[2500],seed[3241],seed[4025],seed[2719],seed[315],seed[3702],seed[1031],seed[3448],seed[1189],seed[3369],seed[3159],seed[3144],seed[3976],seed[3959],seed[3737],seed[1954],seed[1253],seed[3118],seed[3752],seed[2452],seed[1156],seed[1701],seed[2473],seed[191],seed[2174],seed[3772],seed[3523],seed[165],seed[3],seed[2188],seed[1374],seed[2876],seed[3974],seed[3519],seed[3945],seed[2603],seed[2939],seed[3545],seed[912],seed[565],seed[184],seed[1566],seed[1091],seed[2890],seed[1918],seed[1346],seed[1745],seed[3482],seed[2348],seed[3933],seed[3738],seed[2275],seed[1898],seed[2225],seed[667],seed[3092],seed[2612],seed[3193],seed[672],seed[474],seed[1117],seed[830],seed[3023],seed[3967],seed[2061],seed[3416],seed[494],seed[54],seed[3711],seed[3804],seed[1772],seed[1188],seed[2925],seed[2208],seed[1721],seed[3051],seed[3152],seed[3800],seed[2144],seed[1860],seed[2391],seed[3289],seed[1165],seed[3631],seed[289],seed[3769],seed[232],seed[3848],seed[2775],seed[2856],seed[3210],seed[2281],seed[2729],seed[1989],seed[686],seed[605],seed[600],seed[296],seed[706],seed[1514],seed[1029],seed[2744],seed[2148],seed[1221],seed[2336],seed[3376],seed[48],seed[435],seed[179],seed[2232],seed[450],seed[222],seed[2546],seed[3323],seed[3451],seed[1785],seed[895],seed[2987],seed[3420],seed[3763],seed[1248],seed[3546],seed[3319],seed[234],seed[2171],seed[2032],seed[2852],seed[1818],seed[3892],seed[3735],seed[2815],seed[2214],seed[3869],seed[880],seed[293],seed[4049],seed[908],seed[3388],seed[23],seed[193],seed[3398],seed[2367],seed[2785],seed[2062],seed[2832],seed[2875],seed[684],seed[1534],seed[2374],seed[2977],seed[1298],seed[3741],seed[3993],seed[990],seed[2080],seed[2972],seed[3039],seed[1869],seed[3937],seed[722],seed[3133],seed[2313],seed[1862],seed[2924],seed[556],seed[3455],seed[1573],seed[1479],seed[1637],seed[1760],seed[3175],seed[2961],seed[2012],seed[1223],seed[56],seed[2897],seed[2958],seed[141],seed[641],seed[2776],seed[679],seed[3204],seed[2916],seed[1623],seed[624],seed[6],seed[1606],seed[887],seed[2441],seed[2203],seed[491],seed[31],seed[3687],seed[886],seed[118],seed[2695],seed[1369],seed[242],seed[341],seed[2429],seed[736],seed[81],seed[217],seed[2349],seed[285],seed[3947],seed[3064],seed[847],seed[2940],seed[1702],seed[1983],seed[4053],seed[1409],seed[2077],seed[3831],seed[2125],seed[57],seed[2694],seed[1825],seed[1587],seed[3958],seed[905],seed[1469],seed[1145],seed[1146],seed[3254],seed[58],seed[2254],seed[1484],seed[935],seed[625],seed[3872],seed[3243],seed[3704],seed[2150],seed[659],seed[2787],seed[1366],seed[3679],seed[796],seed[1262],seed[3795],seed[1526],seed[3391],seed[2209],seed[2720],seed[1415],seed[3399],seed[2183],seed[909],seed[3893],seed[2094],seed[3557],seed[115],seed[3169],seed[3362],seed[3575],seed[1361],seed[160],seed[3279],seed[2874],seed[1986],seed[1264],seed[2579],seed[4066],seed[542],seed[3748],seed[2172],seed[1037],seed[1889],seed[496],seed[2921],seed[1457],seed[3707],seed[3585],seed[124],seed[2205],seed[778],seed[1905],seed[874],seed[1811],seed[1981],seed[3765],seed[2413],seed[2946],seed[3996],seed[3624],seed[3879],seed[4020],seed[1182],seed[1125],seed[1422],seed[1057],seed[1104],seed[1399],seed[3146],seed[951],seed[236],seed[476],seed[1102],seed[428],seed[3598],seed[1742],seed[2806],seed[2831],seed[1870],seed[2053],seed[2347],seed[871],seed[2202],seed[793],seed[1489],seed[4021],seed[3234],seed[1713],seed[488],seed[3125],seed[3955],seed[3314],seed[2731],seed[2833],seed[2325],seed[3132],seed[2918],seed[2056],seed[287],seed[1666],seed[2492],seed[396],seed[1873],seed[1320],seed[1709],seed[2701],seed[2982],seed[1957],seed[51],seed[824],seed[2434],seed[1080],seed[2189],seed[270],seed[2107],seed[21],seed[692],seed[67],seed[3460],seed[3017],seed[1744],seed[2545],seed[1845],seed[810],seed[1011],seed[2754],seed[527],seed[228],seed[1914],seed[2051],seed[3544],seed[2854],seed[3253],seed[1122],seed[834],seed[462],seed[152],seed[1795],seed[3956],seed[1173],seed[1284],seed[465],seed[1669],seed[1678],seed[3724],seed[3574],seed[3633],seed[812],seed[340],seed[1222],seed[946],seed[2462],seed[3389],seed[2591],seed[660],seed[3621],seed[2634],seed[243],seed[3616],seed[1736],seed[562],seed[1046],seed[3508],seed[2190],seed[117],seed[3662],seed[1071],seed[1302],seed[3517],seed[2532],seed[2409],seed[2200],seed[214],seed[1392],seed[3651],seed[1815],seed[3000],seed[1114],seed[2292],seed[1881],seed[2438],seed[1627],seed[1271],seed[3790],seed[1943],seed[2031],seed[1106],seed[1454],seed[2613],seed[3290],seed[894],seed[1908],seed[3299],seed[101],seed[2238],seed[3541],seed[1228],seed[646],seed[2960],seed[1299],seed[936],seed[32],seed[3353],seed[3818],seed[369],seed[2879],seed[1225],seed[2684],seed[756],seed[1378],seed[311],seed[2377],seed[2375],seed[3529],seed[1580],seed[2446],seed[1564],seed[3918],seed[2196],seed[2396],seed[458],seed[1150],seed[1948],seed[64],seed[1230],seed[962],seed[937],seed[3719],seed[18],seed[2319],seed[2919],seed[2416],seed[602],seed[917],seed[3145],seed[1441],seed[3358],seed[2767],seed[2993],seed[3954],seed[2386],seed[2226],seed[3410],seed[3811],seed[2499],seed[1915],seed[400],seed[3292],seed[3564],seed[3224],seed[1313],seed[3649],seed[2153],seed[1931],seed[913],seed[3718],seed[3059],seed[747],seed[975],seed[2882],seed[3759],seed[1602],seed[3022],seed[1556],seed[901],seed[1509],seed[2649],seed[2311],seed[1432],seed[1330],seed[1730],seed[680],seed[3692],seed[560],seed[3480],seed[3664],seed[1756],seed[2070],seed[2333],seed[3609],seed[3659],seed[212],seed[1413],seed[573],seed[2233],seed[1307],seed[1375],seed[2035],seed[3356],seed[2855],seed[156],seed[1681],seed[1238],seed[4042],seed[1231],seed[3632],seed[2381],seed[2550],seed[2635],seed[3771],seed[3732],seed[467],seed[159],seed[3340],seed[3870],seed[2242],seed[1382],seed[2949],seed[3060],seed[132],seed[441],seed[1644],seed[1612],seed[2025],seed[1407],seed[642],seed[2569],seed[3647],seed[4064],seed[11],seed[2504],seed[1069],seed[1486],seed[3414],seed[2525],seed[2166],seed[1344],seed[2920],seed[2425],seed[3843],seed[1476],seed[3121],seed[1015],seed[1119],seed[3113],seed[2655],seed[38],seed[2024],seed[2294],seed[3478],seed[412],seed[1647],seed[1211],seed[70],seed[526],seed[2942],seed[1471],seed[1343],seed[1993],seed[3345],seed[3819],seed[1097],seed[1021],seed[3932],seed[2727],seed[456],seed[1517],seed[3677],seed[3467],seed[13],seed[1532],seed[700],seed[3646],seed[3239],seed[269],seed[1105],seed[317],seed[561],seed[1690],seed[1028],seed[3231],seed[558],seed[3371],seed[3163],seed[1408],seed[1003],seed[2469],seed[205],seed[3881],seed[1646],seed[4008],seed[1017],seed[2804],seed[2524],seed[1226],seed[1968],seed[2643],seed[1675],seed[202],seed[3427],seed[1095],seed[1662],seed[2857],seed[1595],seed[24],seed[1160],seed[85],seed[885],seed[1495],seed[2605],seed[1970],seed[882],seed[2650],seed[791],seed[3257],seed[2570],seed[889],seed[925],seed[2888],seed[3306],seed[3071],seed[2173],seed[3844],seed[3463],seed[1158],seed[3309],seed[1657],seed[2554],seed[295],seed[1326],seed[2157],seed[334],seed[2165],seed[3046],seed[892],seed[3173],seed[1333],seed[499],seed[1880],seed[3419],seed[279],seed[3461],seed[918],seed[72],seed[3320],seed[3781],seed[931],seed[2991],seed[1635],seed[3225],seed[2320],seed[2585],seed[1782],seed[377],seed[3762],seed[4011],seed[775],seed[3630],seed[4083],seed[2562],seed[1239],seed[3223],seed[2926],seed[701],seed[1244],seed[1072],seed[1208],seed[1490],seed[290],seed[1137],seed[4028],seed[989],seed[1459],seed[3318],seed[1773],seed[53],seed[636],seed[1572],seed[1492],seed[1420],seed[3563],seed[3999],seed[2006],seed[1590],seed[2406],seed[4022],seed[1010],seed[1162],seed[1836],seed[3015],seed[675],seed[3805],seed[508],seed[2820],seed[3502],seed[2783],seed[3250],seed[1498],seed[49],seed[1824],seed[2088],seed[1254],seed[1079],seed[2565],seed[43],seed[699],seed[3526],seed[2072],seed[845],seed[3283],seed[2703],seed[1306],seed[1727],seed[3527],seed[2512],seed[1099],seed[1483],seed[2606],seed[1294],seed[767],seed[4050],seed[1965],seed[997],seed[1296],seed[1448],seed[1466],seed[1205],seed[1309],seed[613],seed[668],seed[1875],seed[691],seed[4069],seed[2089],seed[3591],seed[3981],seed[3982],seed[530],seed[73],seed[1485],seed[3192],seed[1844],seed[162],seed[3165],seed[1329],seed[1741],seed[3683],seed[576],seed[2625],seed[3776],seed[17],seed[3709],seed[1684],seed[1438],seed[1136],seed[1365],seed[1955],seed[622],seed[1118],seed[1243],seed[402],seed[1058],seed[2228],seed[3242],seed[1978],seed[178],seed[2668],seed[3200],seed[911],seed[3890],seed[2706],seed[3571],seed[1397],seed[2536],seed[3150],seed[2461],seed[482],seed[2104],seed[534],seed[2581],seed[4072],seed[2318],seed[2314],seed[1529],seed[3301],seed[1039],seed[868],seed[3127],seed[3528],seed[1376],seed[1679],seed[3422],seed[3579],seed[4038],seed[2989],seed[3106],seed[579],seed[3317],seed[3636],seed[1052],seed[3911],seed[257],seed[1909],seed[853],seed[2661],seed[2795],seed[3876],seed[2432],seed[2139],seed[1446],seed[677],seed[2734],seed[2828],seed[4044],seed[3001],seed[1372],seed[2118],seed[765],seed[254],seed[3619],seed[2930],seed[1683],seed[3815],seed[1694],seed[3382],seed[963],seed[2911],seed[4043],seed[19],seed[2170],seed[1428],seed[1515],seed[3595],seed[861],seed[280],seed[1996],seed[3364],seed[3185],seed[2521],seed[3886],seed[2194],seed[3499],seed[2970],seed[741],seed[2704],seed[571],seed[218],seed[1754],seed[1753],seed[1589],seed[3147],seed[2759],seed[3897],seed[3005],seed[2578],seed[1770],seed[2267],seed[2101],seed[954],seed[2355],seed[2129],seed[1281],seed[2155],seed[688],seed[28],seed[4074],seed[1823],seed[2136],seed[671],seed[1398],seed[1391],seed[1883],seed[2629],seed[717],seed[1591],seed[1184],seed[897],seed[140],seed[1839],seed[627],seed[3614],seed[2866],seed[1135],seed[2867],seed[3026],seed[1194],seed[442],seed[1807],seed[750],seed[3569],seed[1579],seed[1771],seed[1077],seed[2733],seed[238],seed[2475],seed[626],seed[2909],seed[693],seed[2193],seed[2842],seed[3172],seed[3511],seed[548],seed[4060],seed[1703],seed[3442],seed[2711],seed[3908],seed[1009],seed[3164],seed[2191],seed[2531],seed[256],seed[4077],seed[3031],seed[2305],seed[3076],seed[705],seed[942],seed[3884],seed[119],seed[1963],seed[3251],seed[2551],seed[196],seed[2241],seed[3644],seed[1596],seed[888],seed[1363],seed[2906],seed[168],seed[61],seed[944],seed[2738],seed[815],seed[353],seed[490],seed[420],seed[2933],seed[107],seed[1442],seed[3678],seed[3394],seed[209],seed[593],seed[2928],seed[188],seed[1318],seed[3395],seed[3417],seed[2935],seed[2015],seed[3970],seed[998],seed[837],seed[263],seed[799],seed[2580],seed[2162],seed[3612],seed[2732],seed[498],seed[2085],seed[2253],seed[339],seed[1387],seed[2889],seed[1765],seed[1133],seed[2098],seed[2752],seed[923],seed[2127],seed[3313],seed[3434],seed[367],seed[924],seed[323],seed[2788],seed[3122],seed[485],seed[2197],seed[3568],seed[2398],seed[1973],seed[2114],seed[380],seed[3007],seed[2286],seed[3070],seed[1103],seed[740],seed[2519],seed[3975],seed[575],seed[719],seed[2236],seed[780],seed[1600],seed[3924],seed[2100],seed[3255],seed[2250],seed[2664],seed[2937],seed[1604],seed[1935],seed[708],seed[3062],seed[2244],seed[566],seed[1837],seed[1240],seed[1977],seed[1601],seed[1940],seed[3653],seed[698],seed[154],seed[3658],seed[3216],seed[505],seed[729],seed[1452],seed[3035],seed[1658],seed[2862],seed[1123],seed[2681],seed[3774],seed[3274],seed[1171],seed[3003],seed[9],seed[3390],seed[835],seed[981],seed[2686],seed[2677],seed[2608],seed[1138],seed[884],seed[2567],seed[2496],seed[4091],seed[1872],seed[2886],seed[3605],seed[1279],seed[2626],seed[966],seed[3867],seed[3112],seed[3349],seed[2028],seed[2397],seed[2747],seed[587],seed[430],seed[2474],seed[1084],seed[3909],seed[2237],seed[519],seed[3566],seed[2296],seed[100],seed[2383],seed[3377],seed[303],seed[3027],seed[1789],seed[1530],seed[1368],seed[3668],seed[3138],seed[2953],seed[3757],seed[25],seed[2662],seed[3272],seed[1512],seed[305],seed[3428],seed[3550],seed[3657],seed[1491],seed[4058],seed[327],seed[3180],seed[3304],seed[2830],seed[858],seed[960],seed[2627],seed[3565],seed[2248],seed[189],seed[2334],seed[2637],seed[2604],seed[2883],seed[3828],seed[4023],seed[2887],seed[133],seed[343],seed[3931],seed[2354],seed[1013],seed[2530],seed[3114],seed[2628],seed[4095],seed[580],seed[2332],seed[3900],seed[3196],seed[1668],seed[1000],seed[93],seed[1653],seed[1269],seed[45],seed[720],seed[1094],seed[2130],seed[3935],seed[2054],seed[1859],seed[393],seed[1324],seed[1740],seed[3207],seed[1739],seed[4094],seed[2493],seed[3094],seed[2769],seed[2692],seed[1689],seed[298],seed[233],seed[3562],seed[1819],seed[250],seed[2722],seed[103],seed[170],seed[2186],seed[2617],seed[3044],seed[1075],seed[515],seed[985],seed[2063],seed[2638],seed[2086],seed[2274],seed[940],seed[520],seed[4040],seed[3602],seed[1332],seed[1700],seed[2724],seed[2224],seed[1788],seed[1101],seed[3570],seed[2204],seed[2966],seed[3780],seed[3750],seed[3435],seed[545],seed[1331],seed[1256],seed[1038],seed[1947],seed[1073],seed[3174],seed[2278],seed[2756],seed[1733],seed[3663],seed[1886],seed[2428],seed[1074],seed[1801],seed[3220],seed[2824],seed[484],seed[2103],seed[4027],seed[3019],seed[3458],seed[852],seed[1747],seed[2900],seed[2520],seed[866],seed[967],seed[570],seed[1445],seed[900],seed[2528],seed[1502],seed[2690],seed[1018],seed[1803],seed[207],seed[1110],seed[1494],seed[4018],seed[1187],seed[930],seed[811],seed[3934],seed[3135],seed[948],seed[955],seed[1656],seed[3930],seed[142],seed[1799],seed[1798],seed[1991],seed[609],seed[725],seed[2351],seed[451],seed[46],seed[893],seed[2589],seed[3796],seed[1791],seed[3066],seed[1691],seed[3838],seed[3247],seed[1334],seed[974],seed[1643],seed[596],seed[2109],seed[510],seed[559],seed[3342],seed[2652],seed[2050],seed[225],seed[4033],seed[1548],seed[1535],seed[445],seed[3346],seed[1435],seed[1276],seed[820],seed[2300],seed[3149],seed[3847],seed[3643],seed[2517],seed[982],seed[2303],seed[1167],seed[657],seed[3987],seed[1393],seed[1642],seed[2871],seed[4063],seed[2647],seed[1899],seed[2509],seed[199],seed[3871],seed[3964],seed[172],seed[770],seed[739],seed[497],seed[3797],seed[1813],seed[2790],seed[1047],seed[3407],seed[3311],seed[523],seed[1651],seed[3807],seed[589],seed[2584],seed[3661],seed[1624],seed[1323],seed[3885],seed[2751],seed[1796],seed[2914],seed[1060],seed[200],seed[976],seed[3120],seed[2680],seed[732],seed[3977],seed[2247],seed[1107],seed[2648],seed[2936],seed[1050],seed[1923],seed[2192],seed[1603],seed[74],seed[42],seed[486],seed[3782],seed[1019],seed[1421],seed[1885],seed[2199],seed[2586],seed[3137],seed[3904],seed[1115],seed[1149],seed[106],seed[3441],seed[2540],seed[3468],seed[2847],seed[1810],seed[2415],seed[2705],seed[318],seed[2571],seed[2122],seed[346],seed[2400],seed[3720],seed[3214],seed[2757],seed[2894],seed[3827],seed[1381],seed[2152],seed[2252],seed[3115],seed[2548],seed[734],seed[1976],seed[372],seed[16],seed[3922],seed[3655],seed[2723],seed[466],seed[947],seed[619],seed[3091],seed[2384],seed[1834],seed[335],seed[1132],seed[422],seed[1035],seed[447],seed[2380],seed[1168],seed[792],seed[2597],seed[4087],seed[153],seed[516],seed[3509],seed[3852],seed[113],seed[3156],seed[2908],seed[715],seed[87],seed[2913],seed[2881],seed[1628],seed[469],seed[1116],seed[1519],seed[1650],seed[314],seed[1425],seed[1386],seed[2353],seed[763],seed[3012],seed[1664],seed[2147],seed[3963],seed[3587],seed[1577],seed[2800],seed[755],seed[2687],seed[2310],seed[3088],seed[3808],seed[1082],seed[512],seed[4093],seed[1261],seed[1750],seed[1586],seed[584],seed[164],seed[3770],seed[3586],seed[2817],seed[3421],seed[1453],seed[2346],seed[585],seed[2485],seed[760],seed[403],seed[359],seed[1447],seed[2036],seed[2276],seed[3183],seed[2002],seed[2295],seed[4086],seed[1025],seed[2120],seed[551],seed[779],seed[1542],seed[3043],seed[3171],seed[3303],seed[2598],seed[3731],seed[2577],seed[2411],seed[3915],seed[1990],seed[3648],seed[2892],seed[1338],seed[1242],seed[3244],seed[3049],seed[2903],seed[3086],seed[2337],seed[1626],seed[906],seed[2182],seed[653],seed[3433],seed[371],seed[821],seed[55],seed[2742],seed[1195],seed[1636],seed[3676],seed[2113],seed[864],seed[3312],seed[3803],seed[1144],seed[3613],seed[398],seed[4029],seed[2071],seed[4055],seed[210],seed[2027],seed[1516],seed[2359],seed[1578],seed[1051],seed[261],seed[1219],seed[3424],seed[3179],seed[1800],seed[3953],seed[2688],seed[3874],seed[3494],seed[3601],seed[3412],seed[22],seed[768],seed[1549],seed[2312],seed[1894],seed[1067],seed[1555],seed[3045],seed[1615],seed[1599],seed[1109],seed[673],seed[1569],seed[3902],seed[88],seed[532],seed[146],seed[366],seed[221],seed[479],seed[3310],seed[3578],seed[3227],seed[2003],seed[2985],seed[4054],seed[2014],seed[392],seed[814],seed[2670],seed[547],seed[487],seed[489],seed[977],seed[2774],seed[1233],seed[2772],seed[3802],seed[333],seed[1086],seed[360],seed[1098],seed[3308],seed[3073],seed[3627],seed[144],seed[2126],seed[986],seed[2019],seed[1699],seed[2405],seed[1315],seed[408],seed[1697],seed[1980],seed[2097],seed[348],seed[3703],seed[1768],seed[968],seed[3334],seed[3939],seed[3042],seed[2766],seed[3139],seed[2557],seed[1728],seed[2917],seed[1865],seed[3503],seed[3793],seed[2675],seed[1463],seed[1157],seed[1575],seed[2273],seed[1757],seed[1056],seed[255],seed[3286],seed[71],seed[123],seed[2730],seed[929],seed[1449],seed[3277],seed[524],seed[2285],seed[3957],seed[108],seed[3588],seed[1582],seed[150],seed[4046],seed[1288],seed[3457],seed[3691],seed[3926],seed[2878],seed[3866],seed[2301],seed[3929],seed[95],seed[1958],seed[30],seed[223],seed[599],seed[3787],seed[752],seed[2676],seed[2860],seed[3938],seed[3534],seed[2201],seed[62],seed[2042],seed[3298],seed[1561],seed[1474],seed[3829],seed[3197],seed[2588],seed[3498],seed[310],seed[781],seed[2410],seed[3799],seed[1995],seed[3583],seed[39],seed[2389],seed[710],seed[3788],seed[2912],seed[2811],seed[2266],seed[841],seed[2184],seed[2137],seed[2251],seed[397],seed[2083],seed[415],seed[3447],seed[3129],seed[3742],seed[220],seed[3604],seed[216],seed[468],seed[2161],seed[3734],seed[3222],seed[2502],seed[1214],seed[1852],seed[3500],seed[2794],seed[66],seed[1362],seed[3543],seed[1808],seed[643],seed[3756],seed[3328],seed[618],seed[2483],seed[2264],seed[2573],seed[662],seed[1804],seed[2394],seed[1916],seed[3034],seed[1403],seed[338],seed[875],seed[1738],seed[849],seed[1831],seed[3906],seed[3002],seed[586],seed[2582],seed[3488],seed[2243],seed[933],seed[3375],seed[1460],seed[63],seed[1717],seed[854],seed[2671],seed[957],seed[15],seed[3985],seed[773],seed[1439],seed[1994],seed[1988],seed[1890],seed[2282],seed[1111],seed[2073],seed[1410],seed[3794],seed[3952],seed[1436],seed[1054],seed[1966],seed[4034],seed[2735],seed[1351],seed[1673],seed[3998],seed[1480],seed[1280],seed[2636],seed[2302],seed[3916],seed[766],seed[3232],seed[3331],seed[1093],seed[1325],seed[2009],seed[2945],seed[198],seed[370],seed[1934],seed[443],seed[1609],seed[1354],seed[3469],seed[304],seed[336],seed[138],seed[1639],seed[789],seed[416],seed[3491],seed[2641],seed[943],seed[1388],seed[2576],seed[2984],seed[3348],seed[3443],seed[4071],seed[2082],seed[1695],seed[3656],seed[1638],seed[1252],seed[3128],seed[3669],seed[3476],seed[988],seed[2045],seed[1096],seed[631],seed[685],seed[3512],seed[1583],seed[3233],seed[1385],seed[3950],seed[1417],seed[452],seed[128],seed[3010],seed[1175],seed[1780],seed[1776],seed[1164],seed[3905],seed[4079],seed[1864],seed[347],seed[3778],seed[139],seed[682],seed[2457],seed[807],seed[2805],seed[2299],seed[2840],seed[1196],seed[351],seed[1812],seed[2460],seed[111],seed[230],seed[1161],seed[694],seed[2998],seed[2642],seed[3265],seed[116],seed[3567],seed[1998],seed[630],seed[1667],seed[3151],seed[727],seed[301],seed[730],seed[3365],seed[3450],seed[2658],seed[1468],seed[3798],seed[3270],seed[1945],seed[1186],seed[1321],seed[1312],seed[2529],seed[2458],seed[1533],seed[194],seed[3363],seed[829],seed[475],seed[3518],seed[248],seed[405],seed[1204],seed[3625],seed[1210],seed[2240],seed[3177],seed[850],seed[2141],seed[4085],seed[3404],seed[3628],seed[2709],seed[2699],seed[1224],seed[578],seed[3743],seed[3877],seed[1631],seed[564],seed[535],seed[3440],seed[1967],seed[3925],seed[2621],seed[2797],seed[1962],seed[3167],seed[3078],seed[2959],seed[2829],seed[461],seed[3584],seed[2],seed[1303],seed[1500],seed[2623],seed[1607],seed[772],seed[862],seed[2837],seed[3786],seed[1893],seed[2096],seed[928],seed[3611],seed[1622],seed[1250],seed[1551],seed[3104],seed[1982],seed[525],seed[3093],seed[3622],seed[2799],seed[3392],seed[1613],seed[4062],seed[2934],seed[2869],seed[4076],seed[3184],seed[1197],seed[973],seed[3607],seed[246],seed[2466],seed[2872],seed[418],seed[3944],seed[2849],seed[2969],seed[2047],seed[2602],seed[2307],seed[356],seed[1748],seed[1672],seed[1049],seed[3582],seed[2343],seed[3004],seed[3520],seed[4081],seed[3858],seed[1755],seed[1289],seed[978],seed[1121],seed[970],seed[1429],seed[3084],seed[83],seed[1888],seed[1068],seed[2439],seed[2198],seed[337],seed[4089],seed[2269],seed[2372],seed[3266],seed[211],seed[190],seed[3968],seed[714],seed[1680],seed[4092],seed[282],seed[1030],seed[995],seed[539],seed[1652],seed[44],seed[2784],seed[2737],seed[3456],seed[999],seed[2646],seed[1297],seed[536],seed[3332],seed[1353],seed[1632],seed[192],seed[1272],seed[40],seed[3475],seed[2328],seed[4012],seed[1540],seed[2159],seed[2825],seed[3302],seed[4],seed[984],seed[1465],seed[1531],seed[3561],seed[3810],seed[1092],seed[3978],seed[582],seed[1971],seed[2185],seed[477],seed[1112],seed[4045],seed[472],seed[239],seed[473],seed[3832],seed[1383],seed[3733],seed[1305],seed[3134],seed[1896],seed[2339],seed[2067],seed[4004],seed[1024],seed[3912],seed[388],seed[2210],seed[2491],seed[3744],seed[3992],seed[2853],seed[2142],seed[1732],seed[3620],seed[316],seed[2099],seed[3887],seed[1206],seed[2938],seed[746],seed[2683],seed[3271],seed[1707],seed[2000],seed[891],seed[3880],seed[983],seed[650],seed[607],seed[3485],seed[2468],seed[1959],seed[2974],seed[2106],seed[674],seed[2216],seed[1929],seed[938],seed[4001],seed[3402],seed[3888],seed[2124],seed[2904],seed[4059],seed[2566],seed[994],seed[737],seed[3859],seed[3555],seed[3235],seed[608],seed[1611],seed[2119],seed[1621],seed[595],seed[2480],seed[540],seed[2260],seed[3722],seed[1563],seed[563],seed[2081],seed[1126],seed[4088],seed[1659],seed[1268],seed[2345],seed[1283],seed[1719],seed[3357],seed[644],seed[2708],seed[2802],seed[1685],seed[550],seed[1861],seed[2561],seed[3329],seed[3188],seed[1641],seed[2518],seed[439],seed[2026],seed[2331],seed[3535],seed[1040],seed[3530],seed[3385],seed[1558]}),
        .cross_prob(cross_prob),
        .codeword(codeword14),
        .received(received14)
        );
    
    bsc bsc15(
        .clk(clk),
        .reset(reset),
        .seed({seed[603],seed[123],seed[592],seed[851],seed[4074],seed[928],seed[1023],seed[1200],seed[284],seed[1763],seed[566],seed[267],seed[1970],seed[3437],seed[3311],seed[1924],seed[476],seed[3329],seed[2712],seed[2040],seed[526],seed[3334],seed[1001],seed[3335],seed[1408],seed[1523],seed[1945],seed[4093],seed[2339],seed[1895],seed[536],seed[326],seed[887],seed[3034],seed[3885],seed[1885],seed[2805],seed[1343],seed[1144],seed[301],seed[2110],seed[2594],seed[3516],seed[354],seed[1624],seed[3195],seed[1540],seed[72],seed[2421],seed[1340],seed[3116],seed[1549],seed[2385],seed[1626],seed[425],seed[190],seed[1423],seed[2199],seed[1859],seed[1269],seed[1896],seed[1515],seed[2020],seed[3806],seed[4062],seed[1602],seed[1359],seed[938],seed[2679],seed[1092],seed[203],seed[909],seed[1564],seed[2830],seed[482],seed[1159],seed[561],seed[4083],seed[582],seed[2113],seed[389],seed[3048],seed[68],seed[3089],seed[2903],seed[2349],seed[74],seed[2999],seed[3562],seed[3032],seed[3825],seed[1630],seed[2327],seed[744],seed[3850],seed[2375],seed[819],seed[2478],seed[1411],seed[544],seed[4015],seed[2450],seed[3463],seed[1766],seed[2201],seed[455],seed[3384],seed[2939],seed[132],seed[3002],seed[438],seed[1548],seed[4005],seed[1258],seed[3213],seed[2891],seed[699],seed[1636],seed[332],seed[3628],seed[2657],seed[2489],seed[208],seed[325],seed[3888],seed[722],seed[2852],seed[2513],seed[2274],seed[1939],seed[3655],seed[1714],seed[2568],seed[2212],seed[2445],seed[1043],seed[3613],seed[569],seed[2119],seed[4077],seed[1476],seed[554],seed[3193],seed[3889],seed[3391],seed[1202],seed[4043],seed[2610],seed[3462],seed[4054],seed[2018],seed[1058],seed[1036],seed[2543],seed[3596],seed[1000],seed[992],seed[3529],seed[1363],seed[2909],seed[3151],seed[63],seed[3778],seed[3059],seed[3044],seed[1305],seed[1450],seed[3589],seed[1937],seed[172],seed[159],seed[487],seed[1510],seed[899],seed[3107],seed[3421],seed[1122],seed[491],seed[266],seed[2976],seed[146],seed[1274],seed[115],seed[1035],seed[2726],seed[1779],seed[1090],seed[3394],seed[3839],seed[1216],seed[783],seed[2943],seed[3216],seed[3840],seed[2207],seed[486],seed[3123],seed[1625],seed[1740],seed[2680],seed[3261],seed[937],seed[211],seed[2924],seed[794],seed[3077],seed[884],seed[4031],seed[3231],seed[2573],seed[2149],seed[3785],seed[117],seed[1662],seed[3570],seed[3648],seed[2325],seed[3924],seed[4010],seed[1977],seed[2422],seed[1157],seed[2818],seed[3369],seed[3188],seed[3212],seed[1936],seed[743],seed[779],seed[665],seed[2621],seed[3906],seed[657],seed[860],seed[306],seed[112],seed[1729],seed[774],seed[1535],seed[1387],seed[910],seed[2076],seed[2250],seed[413],seed[843],seed[1368],seed[1024],seed[1591],seed[4038],seed[2131],seed[2676],seed[1318],seed[1576],seed[854],seed[3456],seed[1838],seed[2239],seed[3177],seed[3652],seed[2154],seed[1983],seed[639],seed[111],seed[243],seed[629],seed[2273],seed[2300],seed[3321],seed[1691],seed[12],seed[1909],seed[2812],seed[1886],seed[567],seed[1295],seed[350],seed[1586],seed[450],seed[3409],seed[1781],seed[3962],seed[4060],seed[2641],seed[2932],seed[1610],seed[4072],seed[2121],seed[1847],seed[283],seed[3038],seed[3630],seed[189],seed[797],seed[3675],seed[133],seed[1526],seed[2595],seed[1094],seed[2845],seed[2808],seed[1661],seed[2433],seed[2775],seed[648],seed[2703],seed[1638],seed[527],seed[3446],seed[3545],seed[1429],seed[2788],seed[638],seed[3106],seed[1954],seed[898],seed[70],seed[1981],seed[2584],seed[3838],seed[2047],seed[2876],seed[3491],seed[3593],seed[706],seed[18],seed[1210],seed[3954],seed[1427],seed[127],seed[3951],seed[1672],seed[691],seed[749],seed[572],seed[4034],seed[3056],seed[2826],seed[813],seed[1099],seed[1302],seed[249],seed[2384],seed[1064],seed[3362],seed[2918],seed[1809],seed[2326],seed[1645],seed[4088],seed[2078],seed[179],seed[1650],seed[3883],seed[1864],seed[1912],seed[3975],seed[331],seed[109],seed[3173],seed[3257],seed[1021],seed[1456],seed[733],seed[3164],seed[3728],seed[2236],seed[653],seed[2288],seed[2188],seed[2416],seed[1989],seed[3952],seed[836],seed[3587],seed[2534],seed[1826],seed[2254],seed[613],seed[1702],seed[253],seed[120],seed[1979],seed[1760],seed[2564],seed[2637],seed[1160],seed[2900],seed[964],seed[1608],seed[3550],seed[2446],seed[3595],seed[4089],seed[562],seed[3122],seed[3907],seed[186],seed[3285],seed[3015],seed[3070],seed[1491],seed[292],seed[1153],seed[1609],seed[3093],seed[2152],seed[1643],seed[3104],seed[281],seed[40],seed[3941],seed[3606],seed[2752],seed[1335],seed[2803],seed[3688],seed[3897],seed[799],seed[3902],seed[3278],seed[4025],seed[2815],seed[468],seed[1209],seed[2533],seed[1622],seed[215],seed[2605],seed[583],seed[902],seed[1915],seed[1176],seed[1962],seed[1323],seed[2082],seed[3507],seed[859],seed[2695],seed[1304],seed[857],seed[905],seed[3225],seed[2160],seed[1816],seed[1402],seed[472],seed[823],seed[524],seed[2447],seed[3752],seed[980],seed[602],seed[3344],seed[3372],seed[2795],seed[3803],seed[1338],seed[4069],seed[982],seed[251],seed[2869],seed[1765],seed[2650],seed[3694],seed[427],seed[1253],seed[152],seed[3812],seed[1722],seed[3108],seed[1520],seed[311],seed[2569],seed[529],seed[977],seed[3025],seed[1592],seed[636],seed[2180],seed[3232],seed[293],seed[4044],seed[1628],seed[103],seed[1437],seed[3139],seed[2913],seed[2278],seed[2280],seed[3190],seed[875],seed[2111],seed[2714],seed[3567],seed[630],seed[3776],seed[246],seed[1399],seed[3939],seed[4056],seed[1107],seed[556],seed[1453],seed[3672],seed[1517],seed[2243],seed[336],seed[2935],seed[3319],seed[1935],seed[395],seed[2616],seed[3835],seed[1739],seed[3141],seed[1228],seed[563],seed[3283],seed[53],seed[2770],seed[3524],seed[201],seed[57],seed[3660],seed[948],seed[2353],seed[2041],seed[3631],seed[2130],seed[2436],seed[399],seed[1632],seed[2169],seed[280],seed[752],seed[3874],seed[3614],seed[1405],seed[320],seed[2158],seed[145],seed[976],seed[712],seed[1762],seed[3748],seed[1458],seed[2991],seed[2933],seed[3067],seed[3860],seed[1991],seed[2125],seed[1089],seed[3522],seed[3820],seed[2065],seed[36],seed[3789],seed[867],seed[2045],seed[3625],seed[695],seed[1286],seed[2875],seed[1311],seed[698],seed[1529],seed[545],seed[1128],seed[3352],seed[1795],seed[763],seed[116],seed[827],seed[3430],seed[3517],seed[1867],seed[2678],seed[619],seed[3990],seed[999],seed[3185],seed[1412],seed[3417],seed[349],seed[2837],seed[1140],seed[341],seed[3949],seed[2427],seed[3683],seed[50],seed[3144],seed[1310],seed[28],seed[943],seed[2014],seed[3486],seed[892],seed[528],seed[1103],seed[3731],seed[3687],seed[2940],seed[4039],seed[1792],seed[3199],seed[3037],seed[2066],seed[1705],seed[3716],seed[2186],seed[2660],seed[3733],seed[1197],seed[2166],seed[1756],seed[3147],seed[584],seed[1922],seed[2026],seed[3667],seed[1689],seed[2614],seed[3099],seed[1680],seed[49],seed[3588],seed[1759],seed[3821],seed[1439],seed[3057],seed[3330],seed[3131],seed[2737],seed[3503],seed[2997],seed[1347],seed[3314],seed[314],seed[2208],seed[808],seed[1334],seed[1397],seed[3244],seed[1046],seed[500],seed[347],seed[1395],seed[345],seed[1137],seed[3632],seed[2029],seed[371],seed[3339],seed[1240],seed[2490],seed[1623],seed[433],seed[946],seed[3485],seed[1613],seed[392],seed[734],seed[1504],seed[2459],seed[3428],seed[2836],seed[3501],seed[3610],seed[2283],seed[479],seed[3682],seed[1641],seed[2526],seed[2017],seed[2064],seed[4036],seed[3398],seed[2970],seed[3833],seed[1627],seed[2799],seed[1275],seed[3868],seed[304],seed[3434],seed[1278],seed[1279],seed[3348],seed[3512],seed[1522],seed[1749],seed[82],seed[128],seed[3925],seed[3754],seed[929],seed[3980],seed[610],seed[198],seed[1148],seed[1432],seed[2760],seed[2736],seed[969],seed[3496],seed[1919],seed[222],seed[1925],seed[671],seed[2322],seed[418],seed[1357],seed[1553],seed[2256],seed[3324],seed[1300],seed[2484],seed[3247],seed[2746],seed[965],seed[769],seed[2081],seed[1414],seed[1570],seed[1600],seed[2398],seed[3735],seed[1955],seed[4055],seed[3095],seed[1891],seed[2117],seed[512],seed[2864],seed[3197],seed[2059],seed[2221],seed[3921],seed[505],seed[660],seed[1150],seed[4028],seed[192],seed[2839],seed[1670],seed[2509],seed[2898],seed[782],seed[3917],seed[3575],seed[2723],seed[2697],seed[3686],seed[1236],seed[3499],seed[1665],seed[1818],seed[14],seed[2248],seed[3461],seed[1030],seed[3602],seed[2834],seed[3184],seed[259],seed[4012],seed[1131],seed[3282],seed[3965],seed[3742],seed[693],seed[2318],seed[2773],seed[3079],seed[742],seed[221],seed[3206],seed[3872],seed[459],seed[2073],seed[881],seed[2055],seed[380],seed[31],seed[3251],seed[662],seed[3351],seed[3546],seed[805],seed[338],seed[1988],seed[441],seed[1658],seed[791],seed[0],seed[137],seed[1621],seed[560],seed[1114],seed[3011],seed[4051],seed[503],seed[1440],seed[3198],seed[1224],seed[3101],seed[2444],seed[305],seed[1101],seed[1692],seed[815],seed[3645],seed[3696],seed[184],seed[144],seed[2167],seed[1519],seed[2645],seed[3890],seed[3695],seed[3354],seed[3691],seed[2168],seed[2448],seed[3730],seed[3120],seed[3214],seed[1679],seed[3679],seed[2912],seed[3117],seed[907],seed[3412],seed[1882],seed[1356],seed[728],seed[1465],seed[3127],seed[2506],seed[387],seed[1034],seed[2077],seed[2261],seed[1459],seed[2607],seed[853],seed[3337],seed[2298],seed[3192],seed[2463],seed[825],seed[1353],seed[373],seed[2139],seed[2822],seed[3663],seed[1582],seed[183],seed[839],seed[2343],seed[1596],seed[2562],seed[3829],seed[3787],seed[257],seed[2179],seed[3294],seed[2266],seed[2531],seed[3594],seed[3451],seed[844],seed[2783],seed[3792],seed[3992],seed[1798],seed[2833],seed[429],seed[802],seed[1196],seed[188],seed[3920],seed[2311],seed[1797],seed[784],seed[985],seed[3051],seed[9],seed[129],seed[44],seed[1175],seed[2395],seed[69],seed[2219],seed[3904],seed[1799],seed[3218],seed[1085],seed[796],seed[828],seed[1690],seed[118],seed[2787],seed[1676],seed[1881],seed[181],seed[1646],seed[2655],seed[158],seed[2916],seed[2625],seed[3227],seed[3670],seed[1256],seed[3304],seed[3073],seed[166],seed[3571],seed[3264],seed[3256],seed[2690],seed[3714],seed[1449],seed[2380],seed[2608],seed[456],seed[2052],seed[2781],seed[454],seed[272],seed[1289],seed[291],seed[901],seed[3378],seed[3222],seed[2434],seed[2975],seed[2917],seed[3072],seed[962],seed[756],seed[3857],seed[515],seed[3361],seed[1727],seed[3426],seed[1321],seed[3196],seed[2031],seed[3573],seed[1487],seed[1267],seed[2810],seed[3143],seed[1617],seed[2735],seed[212],seed[3438],seed[2780],seed[67],seed[1438],seed[3287],seed[2259],seed[3137],seed[235],seed[3750],seed[1277],seed[1259],seed[2209],seed[2282],seed[3740],seed[581],seed[2871],seed[3183],seed[2617],seed[2520],seed[2128],seed[1127],seed[2499],seed[2216],seed[3822],seed[2418],seed[1095],seed[2],seed[3521],seed[2230],seed[2303],seed[344],seed[3599],seed[4017],seed[3697],seed[2994],seed[3718],seed[1927],seed[1325],seed[3978],seed[861],seed[1163],seed[2681],seed[3246],seed[1180],seed[2659],seed[2571],seed[3404],seed[2269],seed[963],seed[1802],seed[1392],seed[3858],seed[475],seed[1416],seed[1514],seed[740],seed[2959],seed[924],seed[1467],seed[3163],seed[2575],seed[224],seed[1362],seed[504],seed[2794],seed[2604],seed[3782],seed[1785],seed[232],seed[1184],seed[2813],seed[1265],seed[606],seed[4029],seed[403],seed[709],seed[3995],seed[1179],seed[3841],seed[439],seed[2570],seed[2558],seed[3544],seed[838],seed[209],seed[485],seed[1067],seed[1044],seed[1580],seed[1173],seed[1447],seed[3930],seed[3458],seed[1743],seed[918],seed[3482],seed[1499],seed[470],seed[3813],seed[1464],seed[2613],seed[2241],seed[1488],seed[1862],seed[1483],seed[219],seed[2583],seed[1367],seed[3112],seed[1037],seed[353],seed[2831],seed[4006],seed[2858],seed[2175],seed[1509],seed[352],seed[2195],seed[3526],seed[1616],seed[1396],seed[2937],seed[759],seed[1768],seed[240],seed[1100],seed[1551],seed[2860],seed[3725],seed[2357],seed[2027],seed[3909],seed[2290],seed[1307],seed[3415],seed[780],seed[2973],seed[1742],seed[1369],seed[1328],seed[775],seed[758],seed[2423],seed[2734],seed[2574],seed[3064],seed[3910],seed[3474],seed[1857],seed[2846],seed[2715],seed[4094],seed[2372],seed[3489],seed[1109],seed[226],seed[2354],seed[1833],seed[480],seed[227],seed[921],seed[309],seed[2744],seed[787],seed[1422],seed[410],seed[2612],seed[1301],seed[1996],seed[3274],seed[522],seed[3692],seed[3425],seed[1455],seed[1376],seed[2748],seed[33],seed[1139],seed[3024],seed[1492],seed[329],seed[231],seed[3468],seed[1266],seed[711],seed[1250],seed[930],seed[1984],seed[1381],seed[2996],seed[444],seed[3018],seed[3266],seed[2670],seed[587],seed[490],seed[3242],seed[2624],seed[2927],seed[645],seed[2363],seed[1187],seed[4026],seed[754],seed[3781],seed[2165],seed[991],seed[2205],seed[2609],seed[2950],seed[3275],seed[1914],seed[492],seed[1855],seed[3288],seed[1612],seed[661],seed[3542],seed[2386],seed[396],seed[3449],seed[3086],seed[1726],seed[1326],seed[3862],seed[2319],seed[316],seed[4079],seed[550],seed[87],seed[3158],seed[837],seed[1027],seed[3250],seed[2701],seed[2331],seed[187],seed[2244],seed[2656],seed[4087],seed[2694],seed[3230],seed[3745],seed[1571],seed[3423],seed[1640],seed[1585],seed[2778],seed[1388],seed[1642],seed[1629],seed[1928],seed[230],seed[3179],seed[3662],seed[1308],seed[1566],seed[3578],seed[3026],seed[1965],seed[2896],seed[3793],seed[767],seed[2226],seed[1734],seed[2299],seed[3171],seed[2159],seed[1754],seed[2537],seed[2381],seed[981],seed[2136],seed[3472],seed[342],seed[2911],seed[1777],seed[2566],seed[1003],seed[579],seed[631],seed[13],seed[3320],seed[1892],seed[1997],seed[3062],seed[3012],seed[2477],seed[2848],seed[2590],seed[2338],seed[3736],seed[2197],seed[3926],seed[2840],seed[151],seed[2661],seed[3201],seed[2716],seed[3323],seed[2092],seed[30],seed[870],seed[3302],seed[1693],seed[1516],seed[1796],seed[3186],seed[3316],seed[156],seed[1410],seed[1012],seed[3429],seed[202],seed[689],seed[1283],seed[3867],seed[2116],seed[841],seed[2529],seed[612],seed[3022],seed[1011],seed[3987],seed[1557],seed[2948],seed[2790],seed[1126],seed[1942],seed[1306],seed[2265],seed[591],seed[2007],seed[3997],seed[2706],seed[620],seed[2974],seed[564],seed[1312],seed[3142],seed[1195],seed[3654],seed[2630],seed[2036],seed[2494],seed[294],seed[499],seed[2545],seed[2150],seed[1843],seed[3515],seed[1485],seed[2191],seed[2915],seed[2471],seed[2954],seed[3600],seed[3809],seed[961],seed[163],seed[1254],seed[3843],seed[1539],seed[2942],seed[940],seed[1827],seed[96],seed[1025],seed[3871],seed[1226],seed[3895],seed[140],seed[3033],seed[2192],seed[3153],seed[1595],seed[866],seed[1201],seed[3647],seed[3125],seed[3063],seed[3149],seed[1589],seed[2443],seed[2786],seed[481],seed[401],seed[1418],seed[3893],seed[3495],seed[3936],seed[1852],seed[3165],seed[594],seed[416],seed[3615],seed[1717],seed[3050],seed[1911],seed[2341],seed[2741],seed[2144],seed[2161],seed[3295],seed[2765],seed[738],seed[1830],seed[3948],seed[2025],seed[1682],seed[3381],seed[2011],seed[2776],seed[3601],seed[3306],seed[3769],seed[2667],seed[2049],seed[3296],seed[1206],seed[1398],seed[1811],seed[1384],seed[1663],seed[2749],seed[1877],seed[862],seed[2473],seed[2960],seed[2060],seed[973],seed[1614],seed[2557],seed[1272],seed[846],seed[1512],seed[781],seed[2342],seed[3336],seed[4027],seed[258],seed[2229],seed[2387],seed[1169],seed[1124],seed[2989],seed[3317],seed[748],seed[1460],seed[2669],seed[2435],seed[2816],seed[148],seed[3152],seed[3702],seed[1967],seed[2987],seed[960],seed[3475],seed[607],seed[2222],seed[2925],seed[2789],seed[108],seed[1834],seed[3582],seed[2591],seed[3268],seed[1339],seed[351],seed[3592],seed[1309],seed[1284],seed[959],seed[3175],seed[3031],seed[3847],seed[732],seed[2718],seed[3393],seed[1500],seed[4037],seed[3574],seed[2393],seed[3457],seed[2126],seed[2437],seed[2142],seed[2048],seed[372],seed[2091],seed[3366],seed[1031],seed[3103],seed[3454],seed[2177],seed[549],seed[2618],seed[3918],seed[1288],seed[1270],seed[35],seed[967],seed[1652],seed[2333],seed[3756],seed[2348],seed[3309],seed[2185],seed[664],seed[2992],seed[883],seed[1649],seed[3328],seed[900],seed[2072],seed[1771],seed[2184],seed[3642],seed[1587],seed[2213],seed[1873],seed[865],seed[2367],seed[1974],seed[2420],seed[1869],seed[2983],seed[1141],seed[3035],seed[3200],seed[1933],seed[3333],seed[2441],seed[697],seed[1022],seed[2492],seed[1712],seed[2895],seed[3097],seed[2504],seed[2881],seed[674],seed[223],seed[771],seed[2668],seed[3559],seed[1461],seed[2401],seed[713],seed[950],seed[3280],seed[1822],seed[1916],seed[464],seed[2689],seed[4008],seed[3796],seed[1042],seed[1448],seed[3480],seed[1161],seed[414],seed[75],seed[2792],seed[3887],seed[1704],seed[538],seed[3135],seed[92],seed[3611],seed[708],seed[303],seed[1494],seed[3493],seed[58],seed[2408],seed[2552],seed[393],seed[1002],seed[3347],seed[317],seed[2083],seed[2643],seed[3802],seed[3580],seed[2346],seed[1956],seed[1247],seed[3410],seed[1041],seed[3224],seed[2249],seed[2796],seed[1386],seed[995],seed[1478],seed[3661],seed[3955],seed[2947],seed[1923],seed[3643],seed[2855],seed[1181],seed[2811],seed[2798],seed[1725],seed[2977],seed[2090],seed[1102],seed[745],seed[2050],seed[1212],seed[2633],seed[3659],seed[2934],seed[2138],seed[3374],seed[168],seed[3481],seed[1377],seed[904],seed[375],seed[3986],seed[2622],seed[1049],seed[3523],seed[1066],seed[1724],seed[714],seed[1975],seed[3094],seed[2511],seed[2536],seed[457],seed[3259],seed[2291],seed[1213],seed[2647],seed[634],seed[534],seed[3300],seed[1669],seed[795],seed[3514],seed[274],seed[3689],seed[822],seed[1874],seed[1078],seed[210],seed[2003],seed[290],seed[104],seed[376],seed[1020],seed[3401],seed[2698],seed[234],seed[1394],seed[16],seed[390],seed[1477],seed[1987],seed[287],seed[3484],seed[3039],seed[2432],seed[269],seed[942],seed[816],seed[3356],seed[3519],seed[3435],seed[2198],seed[2677],seed[102],seed[1502],seed[1428],seed[2733],seed[1907],seed[2593],seed[2057],seed[3773],seed[86],seed[2100],seed[736],seed[3828],seed[1808],seed[869],seed[1409],seed[3174],seed[2033],seed[2666],seed[1331],seed[3861],seed[3014],seed[1720],seed[3036],seed[176],seed[1425],seed[3360],seed[3269],seed[2938],seed[313],seed[3045],seed[1884],seed[1906],seed[2874],seed[2068],seed[729],seed[3145],seed[2555],seed[2356],seed[886],seed[2133],seed[2944],seed[2337],seed[1993],seed[2865],seed[3617],seed[1647],seed[3439],seed[2493],seed[3864],seed[1770],seed[1684],seed[2360],seed[4033],seed[2646],seed[997],seed[725],seed[237],seed[1863],seed[164],seed[3450],seed[673],seed[25],seed[1593],seed[2464],seed[1918],seed[1681],seed[3935],seed[3923],seed[2628],seed[2549],seed[817],seed[642],seed[465],seed[161],seed[65],seed[3786],seed[2971],seed[2686],seed[2301],seed[2887],seed[333],seed[700],seed[3896],seed[278],seed[1424],seed[2882],seed[1872],seed[1934],seed[2867],seed[1594],seed[3138],seed[3349],seed[3263],seed[718],seed[2129],seed[2215],seed[1578],seed[3898],seed[3364],seed[1075],seed[531],seed[2528],seed[141],seed[1769],seed[383],seed[2252],seed[4068],seed[2482],seed[2019],seed[1940],seed[1832],seed[3541],seed[3946],seed[1010],seed[1950],seed[677],seed[1687],seed[453],seed[3297],seed[340],seed[43],seed[3963],seed[2147],seed[1207],seed[355],seed[1673],seed[2654],seed[3189],seed[3416],seed[1220],seed[1352],seed[2606],seed[2964],seed[3020],seed[1382],seed[1451],seed[3237],seed[3226],seed[3272],seed[2885],seed[2094],seed[134],seed[770],seed[2231],seed[1084],seed[2276],seed[1791],seed[3953],seed[4000],seed[3966],seed[4065],seed[312],seed[2560],seed[248],seed[2889],seed[2310],seed[3815],seed[2980],seed[1055],seed[3508],seed[3299],seed[565],seed[3403],seed[3973],seed[3502],seed[3167],seed[2635],seed[3466],seed[357],seed[3156],seed[296],seed[1846],seed[1840],seed[1132],seed[2819],seed[3612],seed[95],seed[2012],seed[1182],seed[452],seed[1958],seed[100],seed[628],seed[2768],seed[1930],seed[3950],seed[2611],seed[2649],seed[54],seed[2951],seed[3445],seed[1350],seed[510],seed[1198],seed[3724],seed[3794],seed[2880],seed[88],seed[894],seed[1482],seed[1948],seed[1801],seed[702],seed[8],seed[451],seed[2472],seed[2204],seed[692],seed[1960],seed[2945],seed[2268],seed[2228],seed[2620],seed[954],seed[1230],seed[2430],seed[4024],seed[81],seed[588],seed[2227],seed[319],seed[1341],seed[2801],seed[107],seed[1546],seed[1775],seed[1949],seed[658],seed[3157],seed[2350],seed[359],seed[966],seed[3010],seed[245],seed[4059],seed[1992],seed[2108],seed[1573],seed[3510],seed[3389],seed[1841],seed[2523],seed[2114],seed[277],seed[2355],seed[2009],seed[1708],seed[3982],seed[2097],seed[297],seed[914],seed[2894],seed[831],seed[2502],seed[22],seed[97],seed[3098],seed[1471],seed[2352],seed[2086],seed[2955],seed[1233],seed[3365],seed[150],seed[2651],seed[3525],seed[2827],seed[2598],seed[1147],seed[3974],seed[1199],seed[126],seed[3607],seed[3028],seed[1943],seed[2307],seed[1237],seed[3551],seed[1985],seed[1285],seed[182],seed[2403],seed[1214],seed[3845],seed[4092],seed[250],seed[204],seed[2705],seed[1462],seed[3312],seed[2485],seed[2619],seed[3915],seed[1543],seed[1696],seed[647],seed[876],seed[2178],seed[878],seed[366],seed[3999],seed[604],seed[1071],seed[3058],seed[3819],seed[3081],seed[2292],seed[1966],seed[1457],seed[268],seed[2862],seed[2253],seed[580],seed[1844],seed[2683],seed[3598],seed[2340],seed[2998],seed[2242],seed[1648],seed[672],seed[467],seed[3699],seed[1361],seed[1446],seed[3676],seed[2389],seed[1229],seed[3554],seed[3181],seed[3091],seed[3622],seed[3996],seed[2685],seed[788],seed[2507],seed[46],seed[2449],seed[2406],seed[3215],seed[3436],seed[3100],seed[2892],seed[2627],seed[3068],seed[2370],seed[3009],seed[1837],seed[798],seed[2747],seed[3649],seed[2487],seed[1166],seed[398],seed[2731],seed[1978],seed[2275],seed[1401],seed[1655],seed[3236],seed[1825],seed[2196],seed[3976],seed[3041],seed[1496],seed[2551],seed[2272],seed[2383],seed[3090],seed[933],seed[2853],seed[1659],seed[2417],seed[1990],seed[949],seed[270],seed[1611],seed[1635],seed[1372],seed[2601],seed[2402],seed[2724],seed[688],seed[701],seed[814],seed[346],seed[737],seed[3194],seed[2379],seed[1366],seed[1639],seed[1243],seed[2720],seed[680],seed[3658],seed[94],seed[415],seed[2738],seed[1],seed[2688],seed[998],seed[59],seed[2118],seed[986],seed[1248],seed[576],seed[1186],seed[2211],seed[927],seed[3140],seed[1730],seed[2388],seed[739],seed[3082],seed[1231],seed[1653],seed[1081],seed[1105],seed[2329],seed[2907],seed[513],seed[703],seed[1346],seed[3712],seed[1490],seed[557],seed[1737],seed[4022],seed[2691],seed[852],seed[241],seed[2458],seed[2514],seed[1565],seed[2409],seed[2772],seed[1503],seed[3807],seed[2730],seed[2993],seed[1913],seed[2232],seed[2638],seed[945],seed[1773],seed[3539],seed[721],seed[4042],seed[497],seed[2442],seed[3931],seed[2847],seed[3869],seed[365],seed[207],seed[443],seed[821],seed[3397],seed[3770],seed[2106],seed[3407],seed[1820],seed[2439],seed[426],seed[877],seed[3693],seed[1445],seed[682],seed[936],seed[1794],seed[3804],seed[1783],seed[1929],seed[1219],seed[256],seed[3556],seed[2465],seed[681],seed[2956],seed[3238],seed[1544],seed[4003],seed[3638],seed[548],seed[3518],seed[3487],seed[1941],seed[696],seed[2234],seed[2728],seed[411],seed[1545],seed[388],seed[3881],seed[1466],seed[1851],seed[430],seed[167],seed[1061],seed[3],seed[3327],seed[1698],seed[3281],seed[3771],seed[820],seed[21],seed[1480],seed[327],seed[2692],seed[279],seed[2759],seed[1697],seed[2902],seed[1633],seed[521],seed[89],seed[3772],seed[3455],seed[1555],seed[496],seed[3814],seed[3856],seed[449],seed[404],seed[2967],seed[1938],seed[84],seed[3678],seed[2854],seed[85],seed[1415],seed[508],seed[1953],seed[73],seed[142],seed[715],seed[3110],seed[1603],seed[1814],seed[4086],seed[2115],seed[807],seed[2893],seed[911],seed[1865],seed[753],seed[3880],seed[1531],seed[750],seed[1106],seed[3540],seed[76],seed[1959],seed[91],seed[3816],seed[2093],seed[1900],seed[3205],seed[726],seed[934],seed[2016],seed[4058],seed[578],seed[1878],seed[3870],seed[1527],seed[3913],seed[2722],seed[2756],seed[56],seed[4067],seed[2258],seed[147],seed[3380],seed[3779],seed[405],seed[2704],seed[1699],seed[2190],seed[2371],seed[2022],seed[298],seed[2580],seed[3055],seed[1167],seed[2217],seed[3359],seed[328],seed[3969],seed[1508],seed[1706],seed[970],seed[4047],seed[1257],seed[60],seed[381],seed[1518],seed[3007],seed[1009],seed[3768],seed[4073],seed[4045],seed[3467],seed[1108],seed[507],seed[2755],seed[3129],seed[3561],seed[3985],seed[3746],seed[1533],seed[125],seed[3788],seed[667],seed[2286],seed[3853],seed[1736],seed[4070],seed[1174],seed[2453],seed[2474],seed[2921],seed[2260],seed[2067],seed[3379],seed[3154],seed[1964],seed[4048],seed[2470],seed[2366],seed[551],seed[2431],seed[2039],seed[3029],seed[3160],seed[1764],seed[3303],seed[1324],seed[2173],seed[1242],seed[2143],seed[1537],seed[3326],seed[3030],seed[2376],seed[2425],seed[423],seed[3270],seed[1719],seed[3938],seed[1607],seed[539],seed[2302],seed[1619],seed[3075],seed[707],seed[951],seed[2708],seed[618],seed[420],seed[2235],seed[2120],seed[1731],seed[3452],seed[2270],seed[1876],seed[1400],seed[3161],seed[735],seed[1217],seed[979],seed[2127],seed[3916],seed[362],seed[42],seed[1750],seed[2626],seed[1728],seed[1098],seed[2554],seed[2824],seed[3671],seed[2438],seed[3343],seed[773],seed[1403],seed[1858],seed[3558],seed[3836],seed[1282],seed[2214],seed[2218],seed[1436],seed[746],seed[1744],seed[675],seed[1097],seed[29],seed[3584],seed[228],seed[2962],seed[473],seed[1893],seed[1807],seed[760],seed[310],seed[616],seed[3644],seed[121],seed[623],seed[1470],seed[2028],seed[238],seed[1569],seed[3402],seed[407],seed[3492],seed[832],seed[2579],seed[4095],seed[3229],seed[4019],seed[1572],seed[683],seed[3276],seed[1407],seed[2856],seed[590],seed[1281],seed[247],seed[3054],seed[793],seed[27],seed[3134],seed[2396],seed[872],seed[649],seed[1315],seed[2600],seed[932],seed[903],seed[200],seed[2986],seed[3763],seed[2002],seed[3989],seed[2957],seed[1146],seed[1391],seed[3052],seed[3945],seed[2984],seed[1019],seed[687],seed[3709],seed[1417],seed[3624],seed[1047],seed[2546],seed[3826],seed[1441],seed[254],seed[3074],seed[1803],seed[2508],seed[2156],seed[2674],seed[445],seed[1070],seed[178],seed[442],seed[2515],seed[1969],seed[7],seed[1711],seed[422],seed[2246],seed[543],seed[694],seed[428],seed[3548],seed[2561],seed[2483],seed[367],seed[1709],seed[2004],seed[3797],seed[1973],seed[1524],seed[2979],seed[19],seed[199],seed[1303],seed[3879],seed[2978],seed[2255],seed[2793],seed[923],seed[1761],seed[2965],seed[3665],seed[3208],seed[3784],seed[197],seed[3498],seed[379],seed[1443],seed[4057],seed[1133],seed[2308],seed[4085],seed[1618],seed[3531],seed[1668],seed[3605],seed[2632],seed[978],seed[2936],seed[195],seed[3078],seed[1261],seed[2563],seed[1757],seed[1856],seed[840],seed[2577],seed[863],seed[1050],seed[3597],seed[1129],seed[2053],seed[3527],seed[2582],seed[51],seed[3533],seed[2553],seed[3706],seed[3080],seed[1547],seed[1921],seed[3119],seed[261],seed[3656],seed[690],seed[2061],seed[3395],seed[421],seed[3210],seed[540],seed[3774],seed[1980],seed[2105],seed[1378],seed[1143],seed[812],seed[3008],seed[3353],seed[678],seed[3405],seed[1297],seed[2141],seed[2547],seed[2804],seed[2365],seed[2929],seed[1784],seed[1280],seed[3855],seed[2399],seed[1534],seed[1790],seed[2101],seed[656],seed[585],seed[1605],seed[307],seed[322],seed[1014],seed[764],seed[2194],seed[1238],seed[2405],seed[596],seed[3576],seed[3943],seed[1707],seed[171],seed[2306],seed[2132],seed[286],seed[890],seed[3705],seed[3187],seed[3717],seed[384],seed[855],seed[1332],seed[130],seed[1013],seed[1389],seed[52],seed[2429],seed[493],seed[3979],seed[974],seed[3875],seed[3396],seed[1821],seed[3209],seed[633],seed[177],seed[2394],seed[3673],seed[321],seed[3604],seed[3291],seed[1245],seed[893],seed[4035],seed[3536],seed[3345],seed[2522],seed[611],seed[3957],seed[858],seed[2368],seed[1671],seed[1848],seed[1435],seed[2807],seed[1336],seed[2295],seed[1040],seed[397],seed[3873],seed[3202],seed[1191],seed[446],seed[2878],seed[2629],seed[1880],seed[1342],seed[4050],seed[1134],seed[2153],seed[236],seed[2671],seed[3901],seed[3719],seed[1894],seed[2713],seed[2914],seed[2615],seed[3831],seed[3703],seed[2518],seed[553],seed[1452],seed[218],seed[761],seed[983],seed[2838],seed[3087],seed[2001],seed[193],seed[654],seed[3775],seed[3207],seed[1778],seed[285],seed[339],seed[888],seed[1898],seed[3783],seed[3749],seed[3560],seed[1234],seed[2032],seed[2358],seed[1902],seed[1255],seed[1804],seed[2931],seed[2763],seed[830],seed[3377],seed[2411],seed[162],seed[3669],seed[1365],seed[2334],seed[1379],seed[3690],seed[23],seed[988],seed[334],seed[233],seed[3555],seed[3633],seed[2919],seed[2410],seed[3422],seed[2155],seed[3476],seed[3981],seed[2901],seed[48],seed[3668],seed[3367],seed[644],seed[356],seed[2870],seed[2538],seed[1637],seed[776],seed[3228],seed[1971],seed[2104],seed[1317],seed[1004],seed[3811],seed[1944],seed[3998],seed[3292],seed[1138],seed[1287],seed[2099],seed[3385],seed[2098],seed[139],seed[364],seed[2021],seed[1530],seed[1497],seed[3727],seed[3721],seed[1168],seed[1244],seed[1130],seed[2725],seed[1758],seed[2985],seed[2585],seed[3453],seed[3892],seed[2263],seed[3136],seed[1866],seed[806],seed[2497],seed[315],seed[1029],seed[3859],seed[1112],seed[939],seed[3130],seed[1120],seed[2426],seed[3929],seed[1889],seed[1563],seed[913],seed[2884],seed[801],seed[3500],seed[1835],seed[1767],seed[785],seed[2825],seed[595],seed[3162],seed[778],seed[3967],seed[2700],seed[1154],seed[1232],seed[1812],seed[2392],seed[3248],seed[3830],seed[1986],seed[1091],seed[3350],seed[3168],seed[509],seed[3221],seed[2203],seed[2527],seed[3260],seed[532],seed[3220],seed[2440],seed[2843],seed[1561],seed[3027],seed[1532],seed[3239],seed[1904],seed[917],seed[850],seed[2930],seed[947],seed[386],seed[3707],seed[1205],seed[3739],seed[3105],seed[3844],seed[1806],seed[3817],seed[2806],seed[2247],seed[1273],seed[1235],seed[255],seed[824],seed[3085],seed[3651],seed[1276],seed[2897],seed[216],seed[3341],seed[1156],seed[4021],seed[3133],seed[463],seed[2008],seed[2293],seed[2468],seed[206],seed[1579],seed[818],seed[1732],seed[3443],seed[2530],seed[32],seed[3441],seed[1700],seed[915],seed[2777],seed[2135],seed[3933],seed[953],seed[1701],seed[3114],seed[498],seed[3790],seed[2495],seed[2206],seed[157],seed[598],seed[3919],seed[2193],seed[514],seed[165],seed[3734],seed[2157],seed[1223],seed[4023],seed[2817],seed[39],seed[3623],seed[2802],seed[3572],seed[1656],seed[3148],seed[2849],seed[1420],seed[3650],seed[3253],seed[271],seed[1718],seed[358],seed[1963],seed[3286],seed[1604],seed[931],seed[2567],seed[3069],seed[1149],seed[2037],seed[3908],seed[3937],seed[2412],seed[1860],seed[555],seed[4071],seed[2886],seed[2359],seed[1776],seed[2774],seed[3490],seed[1899],seed[2262],seed[1495],seed[3254],seed[3241],seed[1385],seed[2739],seed[2751],seed[1875],seed[2289],seed[502],seed[1871],seed[747],seed[3488],seed[2267],seed[3406],seed[768],seed[1738],seed[1525],seed[3764],seed[3808],seed[1296],seed[3700],seed[1774],seed[1828],seed[289],seed[1383],seed[1327],seed[64],seed[891],seed[78],seed[1716],seed[2102],seed[3370],seed[517],seed[1678],seed[2923],seed[3626],seed[755],seed[676],seed[1033],seed[6],seed[1360],seed[2320],seed[2279],seed[2754],seed[605],seed[2457],seed[2820],seed[2664],seed[3577],seed[3537],seed[2890],seed[484],seed[1513],seed[1017],seed[546],seed[447],seed[1782],seed[265],seed[10],seed[525],seed[717],seed[1789],seed[3191],seed[3528],seed[1810],seed[987],seed[2095],seed[4016],seed[2451],seed[3387],seed[2565],seed[4014],seed[845],seed[2764],seed[3761],seed[2148],seed[1599],seed[3427],seed[1686],seed[2220],seed[751],seed[3262],seed[1861],seed[1155],seed[2758],seed[1073],seed[3569],seed[3905],seed[11],seed[2044],seed[2103],seed[47],seed[864],seed[3180],seed[252],seed[2005],seed[264],seed[3128],seed[3338],seed[3219],seed[3096],seed[3373],seed[3960],seed[993],seed[2559],seed[2369],seed[2982],seed[3922],seed[3066],seed[1710],seed[180],seed[2062],seed[3799],seed[3780],seed[4020],seed[1079],seed[1111],seed[885],seed[1208],seed[1080],seed[2109],seed[3565],seed[93],seed[242],seed[3016],seed[1348],seed[3590],seed[3109],seed[3315],seed[1479],seed[3390],seed[2088],seed[3083],seed[3944],seed[518],seed[573],seed[436],seed[3657],seed[3408],seed[4049],seed[757],seed[632],seed[952],seed[3509],seed[1060],seed[45],seed[110],seed[3150],seed[4063],seed[834],seed[3603],seed[1145],seed[1069],seed[3471],seed[1688],seed[523],seed[3557],seed[811],seed[723],seed[2024],seed[804],seed[1897],seed[2336],seed[2785],seed[1982],seed[3653],seed[124],seed[1723],seed[3400],seed[955],seed[3641],seed[2397],seed[2578],seed[1746],seed[3115],seed[3852],seed[3267],seed[1552],seed[922],seed[3383],seed[136],seed[3616],seed[363],seed[3543],seed[3534],seed[3609],seed[205],seed[1116],seed[2377],seed[1588],seed[1703],seed[975],seed[3701],seed[2210],seed[2035],seed[2762],seed[1442],seed[1473],seed[3447],seed[2013],seed[1575],seed[2652],seed[2480],seed[1121],seed[719],seed[2709],seed[2966],seed[4061],seed[3988],seed[3755],seed[3293],seed[2257],seed[2390],seed[1188],seed[2866],seed[3504],seed[3233],seed[3332],seed[260],seed[2588],seed[3968],seed[1314],seed[3346],seed[2414],seed[2682],seed[488],seed[458],seed[3203],seed[1952],seed[2469],seed[400],seed[637],seed[3310],seed[1463],seed[906],seed[66],seed[2317],seed[494],seed[3621],seed[849],seed[2910],seed[874],seed[727],seed[1606],seed[643],seed[434],seed[668],seed[3704],seed[2673],seed[2112],seed[2501],seed[1651],seed[2745],seed[1074],seed[3563],seed[1337],seed[374],seed[3713],seed[1831],seed[552],seed[3851],seed[1344],seed[3047],seed[2074],seed[1558],seed[1426],seed[3664],seed[1135],seed[2767],seed[1051],seed[1117],seed[3318],seed[1164],seed[330],seed[1489],seed[220],seed[651],seed[1215],seed[1577],seed[406],seed[3473],seed[2455],seed[2475],seed[1032],seed[762],seed[3766],seed[3170],seed[882],seed[324],seed[1125],seed[1511],seed[2750],seed[3411],seed[2122],seed[4030],seed[1358],seed[2452],seed[3903],seed[2510],seed[2850],seed[1076],seed[1045],seed[2535],seed[2642],seed[2640],seed[1054],seed[24],seed[1419],seed[1824],seed[2233],seed[972],seed[99],seed[1330],seed[3738],seed[2539],seed[1674],seed[1354],seed[437],seed[2707],seed[2344],seed[2328],seed[990],seed[1528],seed[2597],seed[38],seed[1747],seed[3715],seed[1292],seed[2648],seed[2503],seed[3759],seed[1088],seed[2592],seed[2189],seed[1193],seed[2174],seed[1241],seed[1486],seed[3970],seed[3023],seed[2952],seed[318],seed[868],seed[2586],seed[1829],seed[4053],seed[1839],seed[3371],seed[2237],seed[394],seed[1252],seed[1068],seed[716],seed[213],seed[1677],seed[3494],seed[1849],seed[1026],seed[3102],seed[3795],seed[1926],seed[956],seed[3666],seed[3591],seed[1995],seed[2085],seed[1375],seed[2345],seed[2466],seed[2162],seed[3866],seed[79],seed[1931],seed[2711],seed[2672],seed[3325],seed[2809],seed[586],seed[2873],seed[2137],seed[2525],seed[2324],seed[1917],seed[2069],seed[2456],seed[2314],seed[1890],seed[3618],seed[3092],seed[368],seed[1316],seed[650],seed[614],seed[2313],seed[2224],seed[1968],seed[469],seed[1190],seed[3640],seed[1887],seed[3399],seed[1264],seed[2861],seed[627],seed[670],seed[460],seed[1634],seed[2800],seed[2572],seed[1222],seed[2462],seed[1225],seed[2717],seed[941],seed[20],seed[2378],seed[3111],seed[3358],seed[2602],seed[273],seed[1946],seed[1431],seed[3538],seed[2419],seed[1836],seed[377],seed[3848],seed[471],seed[3284],seed[2134],seed[570],seed[2023],seed[391],seed[3357],seed[3886],seed[448],seed[1110],seed[786],seed[2599],seed[2264],seed[626],seed[2251],seed[3947],seed[2928],seed[3322],seed[2335],seed[1178],seed[2883],seed[3639],seed[5],seed[3891],seed[879],seed[2187],seed[871],seed[1615],seed[535],seed[1355],seed[61],seed[1787],seed[2908],seed[772],seed[2176],seed[1505],seed[3386],seed[1421],seed[3088],seed[2784],seed[1521],seed[3927],seed[3235],seed[1484],seed[3155],seed[1299],seed[343],seed[1183],seed[3271],seed[2926],seed[2404],seed[2461],seed[1994],seed[3581],seed[2309],seed[2240],seed[615],seed[873],seed[2505],seed[2743],seed[1598],seed[2071],seed[3223],seed[4080],seed[3849],seed[474],seed[1654],seed[1883],seed[154],seed[3732],seed[1583],seed[155],seed[3674],seed[3424],seed[1083],seed[1434],seed[1721],seed[800],seed[1788],seed[378],seed[1903],seed[3777],seed[608],seed[1685],seed[1349],seed[1568],seed[2000],seed[3912],seed[3723],seed[2428],seed[3431],seed[169],seed[2587],seed[2467],seed[1077],seed[810],seed[1329],seed[2476],seed[2863],seed[1374],seed[3132],seed[803],seed[1657],seed[2823],seed[170],seed[1481],seed[1581],seed[369],seed[944],seed[2969],seed[686],seed[173],seed[2146],seed[2990],seed[3301],seed[710],seed[895],seed[2171],seed[4052],seed[1567],seed[3042],seed[114],seed[1028],seed[1239],seed[1062],seed[106],seed[4013],seed[2362],seed[71],seed[1444],seed[1268],seed[2662],seed[3469],seed[295],seed[1142],seed[574],seed[1056],seed[1177],seed[2968],seed[3991],seed[3720],seed[4076],seed[3568],seed[3977],seed[3737],seed[3758],seed[1104],seed[3884],seed[4064],seed[335],seed[288],seed[1507],seed[3388],seed[1320],seed[600],seed[1910],seed[2163],seed[2075],seed[1823],seed[2906],seed[3961],seed[994],seed[537],seed[1291],seed[3076],seed[3124],seed[2972],seed[466],seed[1113],seed[3307],seed[3846],seed[3801],seed[2481],seed[4007],seed[2145],seed[663],seed[2124],seed[3899],seed[3585],seed[1171],seed[3497],seed[501],seed[3553],seed[175],seed[3046],seed[666],seed[2544],seed[3255],seed[880],seed[3635],seed[3722],seed[3204],seed[2512],seed[1805],seed[3375],seed[3084],seed[2170],seed[3636],seed[4090],seed[2486],seed[2548],seed[3940],seed[1694],seed[3277],seed[3532],seed[2719],seed[601],seed[1772],seed[262],seed[3579],seed[1817],seed[2953],seed[3470],seed[1850],seed[519],seed[2323],seed[2151],seed[3854],seed[1072],seed[916],seed[2835],seed[3684],seed[4018],seed[3744],seed[1868],seed[2872],seed[1845],seed[1574],seed[2107],seed[3172],seed[2710],seed[3448],seed[3876],seed[1541],seed[4032],seed[3342],seed[1018],seed[3934],seed[989],seed[1048],seed[1905],seed[1118],seed[3984],seed[724],seed[2183],seed[3432],seed[113],seed[3619],seed[1560],seed[2821],seed[3460],seed[3298],seed[2277],seed[101],seed[3824],seed[3000],seed[3017],seed[3993],seed[1870],seed[3972],seed[2271],seed[3477],seed[4081],seed[1059],seed[2963],seed[2634],seed[847],seed[2687],seed[3392],seed[1998],seed[2415],seed[848],seed[1413],seed[2859],seed[3726],seed[2140],seed[1165],seed[483],seed[1813],seed[935],seed[2988],seed[4066],seed[143],seed[300],seed[1590],seed[3549],seed[2330],seed[1038],seed[1185],seed[2550],seed[589],seed[2769],seed[511],seed[4084],seed[856],seed[646],seed[2532],seed[3520],seed[1584],seed[3440],seed[2382],seed[3005],seed[1380],seed[1536],seed[105],seed[730],seed[896],seed[282],seed[1170],seed[2351],seed[1430],seed[3065],seed[2294],seed[1493],seed[3832],seed[432],seed[1472],seed[361],seed[1390],seed[731],seed[3040],seed[2779],seed[160],seed[2596],seed[2653],seed[83],seed[217],seed[2056],seed[655],seed[1675],seed[2888],seed[174],seed[2413],seed[3118],seed[1119],seed[641],seed[2844],seed[968],seed[1260],seed[3414],seed[370],seed[3583],seed[3878],seed[971],seed[558],seed[2500],seed[777],seed[4],seed[2832],seed[789],seed[2757],seed[2791],seed[3911],seed[1475],seed[3767],seed[766],seed[1468],seed[3680],seed[495],seed[263],seed[1957],seed[3620],seed[417],seed[1664],seed[3837],seed[1364],seed[2842],seed[1096],seed[835],seed[1052],seed[1246],seed[559],seed[3331],seed[122],seed[3478],seed[2516],seed[229],seed[1745],seed[2123],seed[489],seed[419],seed[4075],seed[2905],seed[765],seed[652],seed[2164],seed[2200],seed[3747],seed[1542],seed[2051],seed[3234],seed[897],seed[541],seed[1039],seed[2904],seed[214],seed[2297],seed[194],seed[2766],seed[3159],seed[2364],seed[2517],seed[3760],seed[3800],seed[1433],seed[3060],seed[2042],seed[15],seed[3071],seed[2899],seed[2321],seed[1158],seed[2038],seed[2521],seed[3289],seed[1498],seed[2287],seed[3547],seed[55],seed[3249],seed[1932],seed[3959],seed[2006],seed[1947],seed[1780],seed[3685],seed[2782],seed[3634],seed[2663],seed[3126],seed[2080],seed[3308],seed[3178],seed[2070],seed[3313],seed[302],seed[1227],seed[3827],seed[2828],seed[984],seed[705],seed[2096],seed[244],seed[919],seed[4002],seed[2084],seed[2316],seed[2922],seed[196],seed[3791],seed[2043],seed[547],seed[3513],seed[3608],seed[3290],seed[669],seed[3710],seed[2920],seed[462],seed[17],seed[3535],seed[3176],seed[1005],seed[299],seed[3279],seed[2496],seed[4078],seed[3741],seed[3211],seed[62],seed[1920],seed[912],seed[1660],seed[571],seed[1406],seed[4004],seed[1136],seed[1371],seed[131],seed[2498],seed[3646],seed[431],seed[3243],seed[2058],seed[1601],seed[1901],seed[926],seed[829],seed[4009],seed[2305],seed[2087],seed[3894],seed[958],seed[2540],seed[599],seed[1842],seed[3465],seed[925],seed[2868],seed[2644],seed[225],seed[2581],seed[440],seed[3698],seed[1819],seed[1293],seed[2304],seed[1800],seed[1854],seed[3169],seed[4082],seed[435],seed[3442],seed[98],seed[3419],seed[609],seed[533],seed[593],seed[1715],seed[1393],seed[568],seed[2631],seed[625],seed[908],seed[37],seed[149],seed[2753],seed[3273],seed[3340],seed[1087],seed[1262],seed[1298],seed[3433],seed[3677],seed[2238],seed[1370],seed[842],seed[2639],seed[3865],seed[577],seed[1786],seed[3382],seed[412],seed[275],seed[3505],seed[3900],seed[1501],seed[3265],seed[2407],seed[3413],seed[3363],seed[185],seed[1319],seed[1713],seed[3217],seed[2460],seed[3418],seed[2312],seed[3863],seed[520],seed[2202],seed[1007],seed[809],seed[3708],seed[3971],seed[478],seed[1620],seed[461],seed[3019],seed[575],seed[2841],seed[3765],seed[2015],seed[4001],seed[1469],seed[1015],seed[1151],seed[3810],seed[2675],seed[135],seed[2172],seed[2576],seed[337],seed[2761],seed[1093],seed[1753],seed[506],seed[1879],seed[3627],seed[530],seed[26],seed[138],seed[617],seed[3586],seed[1667],seed[3121],seed[1644],seed[90],seed[408],seed[3166],seed[3003],seed[3805],seed[3994],seed[1597],seed[4091],seed[2851],seed[3258],seed[1082],seed[1815],seed[1351],seed[2603],seed[2636],seed[2797],seed[1562],seed[1194],seed[2079],seed[635],seed[191],seed[2361],seed[622],seed[3355],seed[2721],seed[2696],seed[3061],seed[385],seed[889],seed[1008],seed[3942],seed[704],seed[2740],seed[2941],seed[3566],seed[2089],seed[1115],seed[2285],seed[621],seed[790],seed[516],seed[826],seed[792],seed[2729],seed[3564],seed[833],seed[3245],seed[2857],seed[1908],seed[2374],seed[2223],seed[3743],seed[1559],seed[3182],seed[2054],seed[3753],seed[1853],seed[1016],seed[1972],seed[2046],seed[1631],seed[2225],seed[1333],seed[3757],seed[3013],seed[424],seed[409],seed[1203],seed[1290],seed[1454],seed[2981],seed[2589],seed[2542],seed[2949],seed[1006],seed[1506],seed[3956],seed[1123],seed[3004],seed[1793],seed[34],seed[1666],seed[1204],seed[382],seed[1221],seed[2742],seed[1294],seed[3842],seed[2347],seed[3637],seed[3818],seed[624],seed[3762],seed[2010],seed[1554],seed[119],seed[2281],seed[323],seed[2829],seed[2877],seed[3479],seed[80],seed[1735],seed[1263],seed[1733],seed[3240],seed[3001],seed[3711],seed[741],seed[3729],seed[1550],seed[3958],seed[41],seed[348],seed[276],seed[1752],seed[2034],seed[2958],seed[996],seed[3305],seed[1162],seed[3751],seed[308],seed[1474],seed[1218],seed[920],seed[2702],seed[1755],seed[720],seed[4046],seed[3252],seed[2181],seed[2693],seed[3877],seed[2391],seed[1961],seed[1152],seed[2454],seed[1373],seed[2699],seed[1251],seed[1888],seed[1065],seed[1951],seed[659],seed[3530],seed[3113],seed[2488],seed[1751],seed[685],seed[2332],seed[3798],seed[1976],seed[2479],seed[2296],seed[1086],seed[3049],seed[2684],seed[1556],seed[597],seed[3006],seed[3464],seed[684],seed[1053],seed[3511],seed[3053],seed[1404],seed[2814],seed[3444],seed[3882],seed[542],seed[1189],seed[2623],seed[3834],seed[2727],seed[1313],seed[239],seed[3506],seed[1172],seed[3146],seed[2771],seed[1211],seed[4040],seed[3043],seed[640],seed[1322],seed[2541],seed[2245],seed[2373],seed[77],seed[1192],seed[2491],seed[2424],seed[3983],seed[2995],seed[477],seed[3483],seed[360],seed[679],seed[3914],seed[2879],seed[4041],seed[402],seed[1683],seed[2315],seed[1695],seed[2182],seed[2946],seed[3420],seed[1345],seed[1748],seed[2030],seed[3368],seed[3552],seed[2400],seed[3964],seed[2556],seed[3932],seed[2658],seed[957],seed[2665],seed[3021],seed[3928],seed[4011],seed[3823],seed[3629],seed[1057],seed[1063],seed[3459],seed[2732],seed[1741],seed[153],seed[1538],seed[1271],seed[1999],seed[2063],seed[2961],seed[1249],seed[3376],seed[3681],seed[2524],seed[2519],seed[2284]}),
        .cross_prob(cross_prob),
        .codeword(codeword15),
        .received(received15)
        );
    
    bsc bsc16(
        .clk(clk),
        .reset(reset),
        .seed({seed[1635],seed[1248],seed[3787],seed[2981],seed[3708],seed[1658],seed[331],seed[2234],seed[3108],seed[572],seed[2986],seed[2698],seed[878],seed[2237],seed[2413],seed[375],seed[3458],seed[3375],seed[3565],seed[525],seed[778],seed[2010],seed[136],seed[3235],seed[503],seed[505],seed[2887],seed[3699],seed[1999],seed[377],seed[1526],seed[3019],seed[3343],seed[2770],seed[2160],seed[1362],seed[2650],seed[3276],seed[3230],seed[4066],seed[731],seed[3619],seed[3483],seed[1798],seed[1187],seed[1971],seed[1638],seed[3579],seed[2028],seed[1790],seed[2992],seed[1889],seed[3764],seed[1218],seed[2086],seed[2289],seed[3029],seed[3963],seed[614],seed[1384],seed[56],seed[1239],seed[1927],seed[1315],seed[1996],seed[1656],seed[3988],seed[2186],seed[1757],seed[246],seed[3612],seed[2632],seed[3778],seed[2282],seed[3297],seed[3937],seed[3053],seed[2674],seed[1848],seed[271],seed[452],seed[2714],seed[1690],seed[1486],seed[803],seed[3745],seed[5],seed[3463],seed[1314],seed[2164],seed[3595],seed[283],seed[3114],seed[2032],seed[850],seed[686],seed[3613],seed[3071],seed[120],seed[3581],seed[2097],seed[2260],seed[490],seed[985],seed[3265],seed[711],seed[3119],seed[1318],seed[3357],seed[3869],seed[1069],seed[1832],seed[2124],seed[3540],seed[4067],seed[2216],seed[581],seed[193],seed[119],seed[1223],seed[796],seed[2339],seed[1051],seed[2752],seed[499],seed[388],seed[4087],seed[311],seed[1551],seed[52],seed[1351],seed[588],seed[3913],seed[1493],seed[994],seed[573],seed[2267],seed[1340],seed[1254],seed[4077],seed[223],seed[3634],seed[4094],seed[3130],seed[3487],seed[2795],seed[3608],seed[1843],seed[3720],seed[1725],seed[1302],seed[1027],seed[1091],seed[1780],seed[3317],seed[81],seed[1162],seed[1045],seed[1079],seed[2743],seed[354],seed[1453],seed[2620],seed[1095],seed[862],seed[2584],seed[2964],seed[1370],seed[2570],seed[1772],seed[1730],seed[2358],seed[1577],seed[1781],seed[433],seed[2672],seed[3022],seed[1132],seed[4090],seed[2299],seed[960],seed[1886],seed[2680],seed[172],seed[1936],seed[555],seed[1116],seed[884],seed[2851],seed[1164],seed[1760],seed[607],seed[3982],seed[467],seed[2214],seed[4095],seed[398],seed[1582],seed[2587],seed[4064],seed[3694],seed[501],seed[2198],seed[3045],seed[3942],seed[3006],seed[2611],seed[3650],seed[1066],seed[1192],seed[387],seed[123],seed[1785],seed[86],seed[2499],seed[892],seed[2170],seed[3417],seed[1661],seed[2586],seed[2720],seed[254],seed[84],seed[1673],seed[2852],seed[3460],seed[2573],seed[3295],seed[3548],seed[836],seed[1020],seed[3628],seed[1716],seed[767],seed[3706],seed[2490],seed[2251],seed[882],seed[2244],seed[205],seed[2414],seed[3426],seed[3534],seed[1035],seed[3535],seed[1783],seed[113],seed[1859],seed[1058],seed[3283],seed[845],seed[3233],seed[2205],seed[1731],seed[2196],seed[421],seed[2412],seed[986],seed[2129],seed[2889],seed[1699],seed[1953],seed[2641],seed[45],seed[3657],seed[187],seed[4084],seed[1556],seed[3921],seed[1289],seed[1853],seed[357],seed[2759],seed[510],seed[3396],seed[683],seed[54],seed[126],seed[911],seed[821],seed[1763],seed[2336],seed[832],seed[695],seed[3618],seed[1436],seed[2746],seed[3399],seed[999],seed[1806],seed[3365],seed[3444],seed[2772],seed[905],seed[1010],seed[1256],seed[3394],seed[628],seed[195],seed[2962],seed[3476],seed[2232],seed[1237],seed[780],seed[1378],seed[2163],seed[1086],seed[913],seed[1748],seed[544],seed[828],seed[3892],seed[2043],seed[4009],seed[2295],seed[2566],seed[2017],seed[2554],seed[958],seed[644],seed[1601],seed[275],seed[3563],seed[649],seed[730],seed[2622],seed[1286],seed[2931],seed[3035],seed[3205],seed[1574],seed[3782],seed[346],seed[2471],seed[3146],seed[265],seed[760],seed[1134],seed[1932],seed[1046],seed[988],seed[540],seed[799],seed[917],seed[3829],seed[3267],seed[3600],seed[1458],seed[3739],seed[1398],seed[889],seed[668],seed[1135],seed[3187],seed[3137],seed[2204],seed[276],seed[1878],seed[1594],seed[2423],seed[2215],seed[1048],seed[613],seed[333],seed[2476],seed[3088],seed[3727],seed[923],seed[834],seed[1750],seed[531],seed[1367],seed[3939],seed[1161],seed[1459],seed[2923],seed[2785],seed[3496],seed[975],seed[3896],seed[2046],seed[1296],seed[3559],seed[787],seed[696],seed[2099],seed[1965],seed[2426],seed[2676],seed[2758],seed[497],seed[238],seed[1136],seed[3202],seed[488],seed[1720],seed[2395],seed[79],seed[2877],seed[895],seed[2867],seed[4025],seed[396],seed[1404],seed[3587],seed[2767],seed[2876],seed[1814],seed[1963],seed[3387],seed[3450],seed[3339],seed[2217],seed[3440],seed[2734],seed[1955],seed[3503],seed[473],seed[1677],seed[1073],seed[1882],seed[3799],seed[3314],seed[2303],seed[3725],seed[1924],seed[1609],seed[838],seed[2292],seed[437],seed[2451],seed[1715],seed[179],seed[2769],seed[1964],seed[738],seed[3260],seed[2799],seed[2835],seed[3515],seed[529],seed[125],seed[873],seed[247],seed[2252],seed[3875],seed[1407],seed[763],seed[3853],seed[3076],seed[2357],seed[3116],seed[1726],seed[1316],seed[2559],seed[543],seed[2280],seed[1081],seed[3555],seed[2172],seed[817],seed[3121],seed[347],seed[2970],seed[439],seed[993],seed[3794],seed[1190],seed[2737],seed[1614],seed[941],seed[3354],seed[73],seed[1209],seed[192],seed[2229],seed[3118],seed[826],seed[3907],seed[3574],seed[3656],seed[2858],seed[9],seed[164],seed[3964],seed[2812],seed[3194],seed[3030],seed[1533],seed[2624],seed[422],seed[129],seed[1445],seed[1560],seed[1349],seed[4079],seed[514],seed[4003],seed[3471],seed[368],seed[2527],seed[3768],seed[1007],seed[3277],seed[520],seed[3944],seed[1155],seed[4054],seed[606],seed[1664],seed[761],seed[229],seed[3220],seed[2513],seed[3929],seed[3226],seed[1800],seed[3959],seed[3724],seed[587],seed[1115],seed[4033],seed[1683],seed[1366],seed[3887],seed[3732],seed[1973],seed[4030],seed[3920],seed[1252],seed[719],seed[1185],seed[62],seed[4020],seed[3954],seed[807],seed[3500],seed[105],seed[1053],seed[1562],seed[944],seed[3814],seed[1128],seed[269],seed[2391],seed[2958],seed[3228],seed[815],seed[1692],seed[1172],seed[1326],seed[2219],seed[3897],seed[1666],seed[626],seed[3298],seed[1141],seed[3624],seed[2512],seed[2440],seed[2702],seed[3863],seed[1672],seed[2987],seed[1186],seed[771],seed[2464],seed[1383],seed[2274],seed[380],seed[2265],seed[2226],seed[2128],seed[3854],seed[1849],seed[3900],seed[1280],seed[3777],seed[1842],seed[2177],seed[946],seed[2056],seed[237],seed[3224],seed[1758],seed[3025],seed[487],seed[1345],seed[1625],seed[2115],seed[1472],seed[2757],seed[1344],seed[485],seed[3369],seed[177],seed[535],seed[2338],seed[3512],seed[617],seed[2378],seed[2728],seed[3360],seed[493],seed[1628],seed[3358],seed[3607],seed[457],seed[1338],seed[2488],seed[14],seed[933],seed[3598],seed[1201],seed[3684],seed[2509],seed[2319],seed[635],seed[1586],seed[3451],seed[3181],seed[3752],seed[1468],seed[3304],seed[527],seed[3240],seed[1225],seed[257],seed[1928],seed[3805],seed[1301],seed[4032],seed[1153],seed[1629],seed[2293],seed[964],seed[679],seed[255],seed[4076],seed[3553],seed[1452],seed[2318],seed[227],seed[833],seed[3385],seed[2917],seed[3832],seed[2550],seed[1372],seed[2626],seed[3671],seed[2397],seed[1170],seed[500],seed[2556],seed[1166],seed[1630],seed[848],seed[2606],seed[1513],seed[3625],seed[1102],seed[1159],seed[2246],seed[3957],seed[3253],seed[3986],seed[2079],seed[3946],seed[1126],seed[3893],seed[1967],seed[2685],seed[829],seed[1015],seed[3824],seed[441],seed[3316],seed[1188],seed[3672],seed[3315],seed[1455],seed[1534],seed[2571],seed[75],seed[181],seed[608],seed[2315],seed[1087],seed[1401],seed[3131],seed[2988],seed[2057],seed[1142],seed[2891],seed[1064],seed[2808],seed[1013],seed[3701],seed[2409],seed[2740],seed[1481],seed[218],seed[618],seed[2220],seed[3862],seed[3651],seed[1558],seed[843],seed[3482],seed[656],seed[1580],seed[290],seed[1879],seed[1307],seed[2590],seed[1568],seed[1382],seed[11],seed[4016],seed[2820],seed[224],seed[585],seed[849],seed[1516],seed[3427],seed[2106],seed[3423],seed[1129],seed[3027],seed[3132],seed[1437],seed[3830],seed[3322],seed[2258],seed[3686],seed[4024],seed[1778],seed[2594],seed[26],seed[3643],seed[3207],seed[2257],seed[855],seed[1423],seed[2608],seed[2742],seed[138],seed[330],seed[3580],seed[3851],seed[2083],seed[676],seed[2472],seed[2037],seed[1840],seed[2076],seed[3200],seed[1868],seed[3902],seed[3028],seed[447],seed[394],seed[660],seed[2657],seed[1290],seed[629],seed[2662],seed[3032],seed[1418],seed[270],seed[423],seed[942],seed[1828],seed[1341],seed[1396],seed[3812],seed[2788],seed[1575],seed[1305],seed[2779],seed[2192],seed[689],seed[579],seed[1475],seed[3818],seed[171],seed[2535],seed[3052],seed[2422],seed[2569],seed[2363],seed[2450],seed[1055],seed[2784],seed[3308],seed[2277],seed[2739],seed[3134],seed[2792],seed[1976],seed[2644],seed[3804],seed[4078],seed[3537],seed[2209],seed[3713],seed[1665],seed[3962],seed[1805],seed[2410],seed[463],seed[3871],seed[1706],seed[3721],seed[1520],seed[64],seed[3243],seed[1860],seed[1460],seed[1782],seed[2651],seed[1968],seed[1959],seed[321],seed[1917],seed[2633],seed[2848],seed[3642],seed[1031],seed[4083],seed[36],seed[996],seed[1641],seed[2945],seed[399],seed[2989],seed[3980],seed[442],seed[2883],seed[2369],seed[3860],seed[3161],seed[3345],seed[260],seed[812],seed[720],seed[819],seed[1392],seed[2591],seed[2582],seed[2560],seed[3278],seed[306],seed[2195],seed[2922],seed[3857],seed[1866],seed[918],seed[610],seed[1517],seed[2839],seed[1266],seed[4056],seed[411],seed[557],seed[1264],seed[2558],seed[1913],seed[1844],seed[3926],seed[160],seed[3490],seed[728],seed[3592],seed[2469],seed[2080],seed[2530],seed[340],seed[2806],seed[1737],seed[464],seed[3227],seed[2415],seed[1371],seed[1143],seed[222],seed[3184],seed[2328],seed[1637],seed[1273],seed[847],seed[1532],seed[402],seed[1105],seed[1140],seed[1283],seed[2087],seed[2311],seed[1705],seed[1989],seed[3763],seed[1240],seed[198],seed[2240],seed[1179],seed[870],seed[3178],seed[758],seed[3825],seed[2996],seed[3519],seed[1538],seed[2343],seed[3705],seed[3185],seed[939],seed[496],seed[672],seed[742],seed[1108],seed[1617],seed[1449],seed[153],seed[1678],seed[2640],seed[3311],seed[3372],seed[400],seed[846],seed[777],seed[2718],seed[3941],seed[1009],seed[2661],seed[2896],seed[3293],seed[2747],seed[703],seed[1138],seed[1297],seed[665],seed[1160],seed[363],seed[3556],seed[1242],seed[3631],seed[1738],seed[2437],seed[59],seed[2007],seed[1230],seed[2899],seed[3873],seed[282],seed[943],seed[3401],seed[2932],seed[1040],seed[3326],seed[1462],seed[3649],seed[978],seed[2176],seed[646],seed[2929],seed[2663],seed[1361],seed[3468],seed[391],seed[85],seed[190],seed[2143],seed[2998],seed[997],seed[3397],seed[813],seed[3215],seed[664],seed[2952],seed[3279],seed[3213],seed[3648],seed[3952],seed[3481],seed[511],seed[2646],seed[677],seed[1523],seed[185],seed[2365],seed[3973],seed[2960],seed[699],seed[2392],seed[317],seed[1615],seed[1885],seed[3232],seed[3470],seed[3066],seed[4089],seed[2436],seed[274],seed[2121],seed[2230],seed[3198],seed[3049],seed[981],seed[132],seed[2404],seed[3918],seed[2708],seed[1888],seed[4072],seed[623],seed[1946],seed[2921],seed[66],seed[1415],seed[1691],seed[1529],seed[1986],seed[453],seed[3390],seed[3932],seed[3433],seed[1576],seed[3856],seed[1454],seed[3239],seed[252],seed[1395],seed[1060],seed[2555],seed[3912],seed[2323],seed[1792],seed[4007],seed[3802],seed[3204],seed[995],seed[2713],seed[1113],seed[2879],seed[3211],seed[359],seed[448],seed[1605],seed[823],seed[897],seed[2574],seed[3036],seed[1700],seed[2557],seed[1708],seed[197],seed[3806],seed[558],seed[3521],seed[955],seed[3465],seed[3415],seed[4039],seed[797],seed[2025],seed[147],seed[3009],seed[3575],seed[934],seed[3868],seed[512],seed[1773],seed[1090],seed[4069],seed[2459],seed[2045],seed[2704],seed[559],seed[1646],seed[2701],seed[3425],seed[1648],seed[2592],seed[3325],seed[725],seed[209],seed[1569],seed[292],seed[1542],seed[2071],seed[3095],seed[3928],seed[2690],seed[2968],seed[3165],seed[1123],seed[1310],seed[3400],seed[3557],seed[3828],seed[974],seed[443],seed[3186],seed[2144],seed[1775],seed[2859],seed[1680],seed[2589],seed[3916],seed[1825],seed[1890],seed[1306],seed[3743],seed[984],seed[586],seed[3518],seed[876],seed[2073],seed[1385],seed[3176],seed[2107],seed[3827],seed[1815],seed[2145],seed[41],seed[1549],seed[1626],seed[2496],seed[1983],seed[4037],seed[3590],seed[2110],seed[582],seed[1940],seed[2673],seed[3632],seed[3622],seed[1279],seed[3287],seed[2473],seed[1444],seed[2810],seed[3193],seed[1198],seed[1098],seed[3975],seed[701],seed[2201],seed[602],seed[2432],seed[3418],seed[2354],seed[1016],seed[2683],seed[2818],seed[2278],seed[3138],seed[1537],seed[3381],seed[1883],seed[1813],seed[899],seed[3785],seed[998],seed[407],seed[2925],seed[1528],seed[3229],seed[2732],seed[80],seed[810],seed[2462],seed[1085],seed[861],seed[3620],seed[783],seed[1573],seed[1291],seed[2390],seed[630],seed[970],seed[3175],seed[3145],seed[2006],seed[888],seed[2933],seed[1590],seed[1078],seed[3439],seed[2327],seed[1911],seed[3583],seed[1751],seed[1490],seed[1662],seed[1521],seed[3728],seed[72],seed[502],seed[343],seed[2030],seed[1104],seed[47],seed[2763],seed[1717],seed[1689],seed[2340],seed[2572],seed[2285],seed[1793],seed[1922],seed[1564],seed[1446],seed[2712],seed[908],seed[3577],seed[2607],seed[118],seed[371],seed[281],seed[2817],seed[2865],seed[416],seed[2691],seed[1895],seed[3221],seed[2502],seed[3610],seed[1548],seed[3864],seed[325],seed[2184],seed[616],seed[1695],seed[710],seed[3442],seed[2537],seed[1281],seed[4010],seed[2202],seed[3816],seed[1795],seed[2719],seed[2168],seed[764],seed[2609],seed[3726],seed[1624],seed[1912],seed[355],seed[980],seed[251],seed[1410],seed[2872],seed[2565],seed[662],seed[621],seed[1246],seed[3323],seed[1313],seed[3978],seed[1257],seed[3850],seed[3955],seed[174],seed[294],seed[605],seed[3740],seed[1364],seed[3395],seed[3309],seed[1175],seed[2910],seed[3508],seed[3710],seed[3709],seed[3301],seed[1325],seed[3539],seed[2302],seed[4],seed[2181],seed[3270],seed[2048],seed[576],seed[4045],seed[53],seed[207],seed[3582],seed[2297],seed[563],seed[781],seed[3344],seed[979],seed[2016],seed[3231],seed[87],seed[948],seed[2012],seed[320],seed[2829],seed[1740],seed[1707],seed[4029],seed[1334],seed[2652],seed[3303],seed[83],seed[2372],seed[1687],seed[1839],seed[1150],seed[454],seed[1319],seed[3330],seed[762],seed[3754],seed[465],seed[2900],seed[2744],seed[3822],seed[2194],seed[184],seed[2489],seed[3685],seed[2705],seed[3536],seed[2875],seed[2287],seed[3691],seed[3605],seed[1328],seed[1583],seed[1921],seed[1089],seed[3441],seed[3434],seed[250],seed[1704],seed[1514],seed[2250],seed[1933],seed[740],seed[3562],seed[1835],seed[0],seed[3288],seed[3089],seed[1269],seed[2005],seed[176],seed[2729],seed[298],seed[713],seed[3674],seed[792],seed[3333],seed[322],seed[3588],seed[3275],seed[2162],seed[3180],seed[3000],seed[2627],seed[1919],seed[611],seed[2174],seed[3696],seed[1251],seed[4012],seed[1623],seed[2508],seed[3846],seed[3569],seed[2070],seed[2088],seed[1434],seed[2157],seed[1891],seed[300],seed[3561],seed[519],seed[428],seed[2974],seed[2761],seed[3596],seed[1465],seed[2724],seed[3750],seed[2826],seed[2183],seed[1747],seed[2361],seed[3],seed[384],seed[358],seed[432],seed[1125],seed[3210],seed[1610],seed[1375],seed[2382],seed[1612],seed[3452],seed[2679],seed[3190],seed[1387],seed[3773],seed[580],seed[3578],seed[1097],seed[3981],seed[2881],seed[312],seed[2843],seed[914],seed[2134],seed[1299],seed[2261],seed[1650],seed[1771],seed[3905],seed[3154],seed[989],seed[2091],seed[734],seed[3015],seed[2044],seed[702],seed[1915],seed[2453],seed[3256],seed[2228],seed[173],seed[6],seed[1600],seed[2693],seed[1808],seed[1212],seed[291],seed[4026],seed[178],seed[3718],seed[750],seed[2773],seed[1850],seed[309],seed[3044],seed[3621],seed[134],seed[263],seed[3192],seed[121],seed[97],seed[264],seed[1694],seed[3408],seed[2098],seed[3584],seed[3055],seed[2478],seed[2920],seed[2643],seed[33],seed[2275],seed[1106],seed[2135],seed[2367],seed[3173],seed[2903],seed[3516],seed[612],seed[2018],seed[124],seed[3447],seed[338],seed[2101],seed[652],seed[1033],seed[2094],seed[1036],seed[1743],seed[1137],seed[3693],seed[2222],seed[1011],seed[3938],seed[1670],seed[1380],seed[3550],seed[3477],seed[1987],seed[3765],seed[2360],seed[2428],seed[2002],seed[953],seed[3082],seed[2616],seed[3646],seed[1505],seed[2790],seed[3532],seed[2371],seed[1916],seed[3286],seed[2211],seed[2778],seed[3876],seed[418],seed[2435],seed[2465],seed[3993],seed[739],seed[1755],seed[3925],seed[2575],seed[2114],seed[504],seed[1711],seed[756],seed[1768],seed[2189],seed[3453],seed[25],seed[2534],seed[2515],seed[1535],seed[2653],seed[1145],seed[3046],seed[2975],seed[1061],seed[3112],seed[3072],seed[726],seed[2544],seed[3527],seed[2716],seed[1657],seed[765],seed[1466],seed[3927],seed[1093],seed[1567],seed[383],seed[2993],seed[1205],seed[2380],seed[3206],seed[3282],seed[2449],seed[492],seed[2431],seed[356],seed[1496],seed[3554],seed[372],seed[3617],seed[2288],seed[2433],seed[1381],seed[189],seed[522],seed[3247],seed[3826],seed[2581],seed[2617],seed[1647],seed[2904],seed[150],seed[151],seed[1679],seed[1447],seed[1732],seed[1259],seed[3086],seed[494],seed[3012],seed[539],seed[1881],seed[3241],seed[2748],seed[3337],seed[794],seed[3681],seed[716],seed[655],seed[2760],seed[4014],seed[2480],seed[589],seed[3122],seed[3169],seed[1030],seed[1443],seed[2294],seed[3890],seed[2182],seed[3984],seed[650],seed[3786],seed[3329],seed[2798],seed[2520],seed[1676],seed[2350],seed[2103],seed[2347],seed[3371],seed[4086],seed[2601],seed[1063],seed[1482],seed[2501],seed[2169],seed[455],seed[3769],seed[2655],seed[231],seed[2753],seed[3968],seed[484],seed[951],seed[2786],seed[546],seed[3074],seed[4046],seed[2159],seed[459],seed[566],seed[2377],seed[3430],seed[3711],seed[2486],seed[395],seed[155],seed[3811],seed[2063],seed[1993],seed[3429],seed[68],seed[1037],seed[1285],seed[3910],seed[1471],seed[2963],seed[140],seed[145],seed[3081],seed[1620],seed[2782],seed[3380],seed[2949],seed[789],seed[2504],seed[406],seed[95],seed[3140],seed[775],seed[288],seed[1148],seed[1803],seed[3623],seed[568],seed[1884],seed[2972],seed[2061],seed[2855],seed[3498],seed[1207],seed[2514],seed[1429],seed[2816],seed[2831],seed[1876],seed[2495],seed[2364],seed[2938],seed[74],seed[601],seed[1421],seed[3393],seed[596],seed[3179],seed[1831],seed[4013],seed[1962],seed[3652],seed[3378],seed[1602],seed[1473],seed[1502],seed[688],seed[1425],seed[1109],seed[2600],seed[1960],seed[749],seed[2588],seed[35],seed[3790],seed[722],seed[3334],seed[3741],seed[2510],seed[3940],seed[3064],seed[2888],seed[1497],seed[506],seed[1177],seed[2916],seed[272],seed[2402],seed[3174],seed[909],seed[1863],seed[1117],seed[89],seed[3057],seed[1920],seed[3070],seed[1197],seed[1952],seed[1184],seed[285],seed[3915],seed[1599],seed[1287],seed[2541],seed[3586],seed[793],seed[71],seed[382],seed[2847],seed[1833],seed[1943],seed[3712],seed[2188],seed[3560],seed[201],seed[3300],seed[1193],seed[3061],seed[746],seed[410],seed[415],seed[2411],seed[1320],seed[1561],seed[2796],seed[3966],seed[1898],seed[4038],seed[133],seed[2154],seed[3110],seed[2055],seed[3100],seed[91],seed[213],seed[2854],seed[65],seed[3788],seed[3488],seed[1120],seed[1413],seed[2730],seed[1552],seed[1167],seed[3517],seed[1288],seed[361],seed[3636],seed[654],seed[390],seed[3819],seed[1622],seed[2109],seed[1801],seed[3217],seed[3789],seed[1820],seed[2850],seed[1660],seed[1713],seed[16],seed[3435],seed[600],seed[3336],seed[348],seed[2000],seed[3965],seed[2457],seed[217],seed[2379],seed[1356],seed[1448],seed[2393],seed[3250],seed[1937],seed[1216],seed[2036],seed[1788],seed[426],seed[1270],seed[339],seed[2108],seed[2003],seed[2642],seed[4088],seed[4055],seed[3058],seed[2243],seed[3328],seed[2648],seed[2985],seed[1871],seed[2546],seed[3269],seed[3771],seed[2033],seed[3775],seed[3678],seed[865],seed[3109],seed[2112],seed[3416],seed[3813],seed[1598],seed[2286],seed[2042],seed[2678],seed[3382],seed[3263],seed[867],seed[2041],seed[1337],seed[161],seed[1753],seed[130],seed[2551],seed[3364],seed[2474],seed[3424],seed[2466],seed[1817],seed[2381],seed[1094],seed[3376],seed[3107],seed[3411],seed[801],seed[592],seed[1227],seed[2756],seed[881],seed[2139],seed[3502],seed[144],seed[2349],seed[1154],seed[2305],seed[859],seed[3274],seed[1034],seed[3048],seed[477],seed[3523],seed[3341],seed[2062],seed[634],seed[1202],seed[2579],seed[550],seed[3351],seed[3606],seed[732],seed[1746],seed[214],seed[1477],seed[3974],seed[4031],seed[2346],seed[864],seed[3128],seed[2687],seed[3983],seed[2629],seed[1234],seed[1304],seed[643],seed[2482],seed[2997],seed[860],seed[903],seed[77],seed[4047],seed[2445],seed[374],seed[169],seed[2442],seed[2052],seed[3105],seed[3037],seed[3919],seed[1492],seed[837],seed[1530],seed[1544],seed[3111],seed[3914],seed[1054],seed[3356],seed[1335],seed[2863],seed[3246],seed[3703],seed[2539],seed[2040],seed[3770],seed[1830],seed[3970],seed[2545],seed[305],seed[2038],seed[2383],seed[1565],seed[715],seed[329],seed[1988],seed[163],seed[2707],seed[1938],seed[3238],seed[2291],seed[32],seed[3747],seed[1906],seed[27],seed[2241],seed[2264],seed[670],seed[1893],seed[3492],seed[168],seed[2185],seed[1480],seed[3059],seed[3366],seed[232],seed[1494],seed[2549],seed[2621],seed[1461],seed[239],seed[751],seed[532],seed[3189],seed[690],seed[1697],seed[717],seed[1518],seed[2517],seed[4063],seed[3735],seed[827],seed[904],seed[3342],seed[444],seed[2425],seed[3249],seed[3697],seed[3865],seed[3318],seed[3626],seed[2930],seed[1762],seed[1639],seed[1284],seed[627],seed[2822],seed[3023],seed[3729],seed[3063],seed[647],seed[542],seed[2647],seed[1408],seed[2446],seed[2950],seed[2585],seed[324],seed[3151],seed[795],seed[2577],seed[2253],seed[491],seed[2388],seed[3248],seed[3738],seed[2825],seed[929],seed[4035],seed[2834],seed[167],seed[1634],seed[1438],seed[2254],seed[2543],seed[1004],seed[2861],seed[127],seed[3704],seed[645],seed[381],seed[3234],seed[2866],seed[2179],seed[3486],seed[2353],seed[3414],seed[1228],seed[2856],seed[1232],seed[3080],seed[2193],seed[641],seed[370],seed[3043],seed[3670],seed[3664],seed[4091],seed[661],seed[2604],seed[874],seed[1826],seed[822],seed[1277],seed[15],seed[1804],seed[1642],seed[1651],seed[157],seed[435],seed[3493],seed[1539],seed[2213],seed[3142],seed[3667],seed[620],seed[2065],seed[755],seed[3011],seed[2631],seed[2765],seed[533],seed[2366],seed[293],seed[3855],seed[1742],seed[2078],seed[1017],seed[3753],seed[1439],seed[2635],seed[1770],seed[2406],seed[413],seed[2939],seed[3969],seed[3067],seed[456],seed[3541],seed[1139],seed[3075],seed[685],seed[3715],seed[1794],seed[536],seed[3096],seed[2552],seed[785],seed[3117],seed[1261],seed[2148],seed[2419],seed[1718],seed[3679],seed[2967],seed[940],seed[2871],seed[651],seed[2845],seed[2484],seed[1873],seed[1221],seed[2180],seed[3604],seed[830],seed[1243],seed[3707],seed[1767],seed[3630],seed[2598],seed[1531],seed[2105],seed[475],seed[2892],seed[707],seed[2069],seed[462],seed[2966],seed[2731],seed[952],seed[1945],seed[3756],seed[2942],seed[1616],seed[2941],seed[3934],seed[2004],seed[3682],seed[3861],seed[741],seed[1667],seed[13],seed[2092],seed[7],seed[2522],seed[1379],seed[624],seed[341],seed[3195],seed[335],seed[2421],seed[2191],seed[262],seed[244],seed[3525],seed[1925],seed[959],seed[3445],seed[342],seed[2399],seed[1816],seed[2233],seed[3284],seed[3392],seed[615],seed[2727],seed[3047],seed[420],seed[637],seed[1595],seed[2959],seed[3412],seed[1350],seed[3148],seed[1961],seed[2138],seed[2533],seed[1038],seed[947],seed[1183],seed[267],seed[2983],seed[3638],seed[3666],seed[1607],seed[191],seed[3877],seed[1572],seed[2123],seed[2256],seed[3759],seed[286],seed[2531],seed[1321],seed[3324],seed[3923],seed[1099],seed[3079],seed[3144],seed[3362],seed[2971],seed[438],seed[3979],seed[3398],seed[3662],seed[852],seed[2368],seed[737],seed[1969],seed[364],seed[1649],seed[2085],seed[574],seed[3888],seed[991],seed[820],seed[1426],seed[1511],seed[636],seed[774],seed[2334],seed[3355],seed[3884],seed[3348],seed[591],seed[1908],seed[2218],seed[3641],seed[1579],seed[3428],seed[2807],seed[352],seed[2681],seed[928],seed[2460],seed[3616],seed[1047],seed[3335],seed[3281],seed[2776],seed[3251],seed[1698],seed[3242],seed[48],seed[334],seed[3403],seed[2401],seed[3208],seed[609],seed[102],seed[2141],seed[389],seed[4036],seed[2862],seed[3083],seed[1627],seed[2783],seed[1399],seed[1174],seed[2583],seed[3528],seed[3924],seed[3901],seed[2269],seed[1684],seed[1734],seed[3084],seed[3489],seed[2630],seed[2122],seed[3796],seed[1841],seed[2936],seed[3338],seed[307],seed[3219],seed[3717],seed[759],seed[863],seed[1491],seed[109],seed[773],seed[2394],seed[2529],seed[2605],seed[1057],seed[570],seed[3160],seed[4041],seed[3222],seed[2692],seed[1929],seed[3167],seed[2781],seed[2578],seed[78],seed[2898],seed[2658],seed[412],seed[2456],seed[3762],seed[2821],seed[2519],seed[1702],seed[3820],seed[2645],seed[3257],seed[3730],seed[373],seed[3158],seed[3254],seed[508],seed[898],seed[3102],seed[297],seed[3010],seed[3272],seed[2787],seed[2084],seed[1709],seed[3629],seed[3368],seed[2116],seed[1092],seed[104],seed[3858],seed[631],seed[1268],seed[3766],seed[2722],seed[806],seed[1008],seed[2072],seed[57],seed[3018],seed[2666],seed[976],seed[1581],seed[2498],seed[1724],seed[3698],seed[1478],seed[598],seed[1838],seed[1176],seed[2823],seed[3669],seed[3472],seed[2173],seed[3776],seed[2344],seed[2384],seed[1896],seed[2800],seed[2766],seed[107],seed[2842],seed[2444],seed[3835],seed[927],seed[3410],seed[234],seed[2161],seed[1352],seed[3683],seed[1653],seed[745],seed[2326],seed[1430],seed[3021],seed[551],seed[3882],seed[3842],seed[3040],seed[887],seed[2126],seed[3880],seed[2373],seed[957],seed[2166],seed[1631],seed[4050],seed[809],seed[1809],seed[2492],seed[3947],seed[1376],seed[2567],seed[2470],seed[3594],seed[2111],seed[1741],seed[1411],seed[3172],seed[642],seed[3259],seed[2307],seed[1854],seed[1433],seed[3599],seed[1072],seed[1118],seed[367],seed[204],seed[1181],seed[790],seed[961],seed[1857],seed[3639],seed[965],seed[2723],seed[1278],seed[916],seed[2158],seed[886],seed[680],seed[240],seed[3404],seed[727],seed[3719],seed[2049],seed[2019],seed[1640],seed[2526],seed[779],seed[3961],seed[110],seed[4015],seed[196],seed[2247],seed[1686],seed[901],seed[4059],seed[2420],seed[2654],seed[301],seed[3383],seed[1956],seed[1173],seed[2483],seed[1761],seed[3113],seed[2832],seed[1931],seed[135],seed[2726],seed[203],seed[3386],seed[405],seed[296],seed[2775],seed[202],seed[1000],seed[128],seed[816],seed[1019],seed[2156],seed[1942],seed[414],seed[2479],seed[1180],seed[1597],seed[2675],seed[597],seed[1984],seed[2901],seed[474],seed[1133],seed[2638],seed[1059],seed[3654],seed[3520],seed[2375],seed[982],seed[137],seed[648],seed[3972],seed[2133],seed[1103],seed[2427],seed[149],seed[480],seed[3702],seed[2564],seed[2880],seed[2669],seed[851],seed[1618],seed[885],seed[386],seed[1570],seed[3748],seed[575],seed[1654],seed[1],seed[76],seed[360],seed[1902],seed[983],seed[4040],seed[3252],seed[378],seed[2059],seed[1926],seed[3737],seed[883],seed[3791],seed[1671],seed[1112],seed[3746],seed[1463],seed[1789],seed[2870],seed[1327],seed[3157],seed[2245],seed[4071],seed[2095],seed[1990],seed[924],seed[2697],seed[736],seed[55],seed[2505],seed[2058],seed[2794],seed[4018],seed[38],seed[673],seed[1200],seed[3546],seed[962],seed[34],seed[1258],seed[3558],seed[561],seed[3547],seed[3817],seed[2325],seed[2497],seed[4043],seed[450],seed[1519],seed[3191],seed[2200],seed[1723],seed[4053],seed[3031],seed[2322],seed[3307],seed[289],seed[1483],seed[2677],seed[3377],seed[43],seed[1076],seed[1196],seed[3120],seed[2239],seed[1331],seed[920],seed[3094],seed[2494],seed[593],seed[2503],seed[3742],seed[249],seed[931],seed[3576],seed[2793],seed[17],seed[1571],seed[3511],seed[3182],seed[1068],seed[2352],seed[2153],seed[2175],seed[3352],seed[1359],seed[2370],seed[4068],seed[4073],seed[1217],seed[1414],seed[2255],seed[2400],seed[2836],seed[709],seed[2348],seed[1507],seed[2356],seed[1923],seed[98],seed[1424],seed[2755],seed[1712],seed[1824],seed[3268],seed[1336],seed[3155],seed[4042],seed[3522],seed[4070],seed[2809],seed[528],seed[287],seed[2523],seed[930],seed[268],seed[3544],seed[800],seed[182],seed[1901],seed[2894],seed[2837],seed[3843],seed[3834],seed[1547],seed[2500],seed[1213],seed[2281],seed[2750],seed[1124],seed[3197],seed[2090],seed[1071],seed[228],seed[3953],seed[714],seed[2946],seed[3609],seed[3209],seed[788],seed[1950],seed[708],seed[2634],seed[482],seed[1157],seed[2104],seed[2853],seed[2660],seed[1353],seed[1215],seed[3319],seed[2051],seed[3614],seed[1644],seed[967],seed[233],seed[1122],seed[1752],seed[108],seed[1948],seed[3676],seed[1796],seed[3585],seed[3551],seed[3042],seed[3513],seed[3722],seed[362],seed[2548],seed[1722],seed[1769],seed[2403],seed[3466],seed[401],seed[115],seed[1158],seed[3549],seed[1119],seed[638],seed[22],seed[1163],seed[3886],seed[154],seed[1342],seed[1836],seed[1080],seed[3236],seed[1373],seed[3680],seed[3781],seed[1765],seed[2113],seed[2602],seed[2331],seed[3419],seed[3744],seed[4017],seed[1088],seed[1100],seed[67],seed[3420],seed[2542],seed[910],seed[2387],seed[2074],seed[2994],seed[1470],seed[2840],seed[1823],seed[3695],seed[3971],seed[1500],seed[2487],seed[1348],seed[1169],seed[857],seed[3005],seed[1555],seed[3087],seed[142],seed[1479],seed[3529],seed[3506],seed[1435],seed[1220],seed[906],seed[4057],seed[345],seed[4052],seed[2454],seed[3056],seed[554],seed[769],seed[782],seed[2937],seed[3815],seed[3153],seed[3407],seed[3289],seed[972],seed[3150],seed[3542],seed[2385],seed[3573],seed[2026],seed[2689],seed[3361],seed[1365],seed[3690],seed[772],seed[2736],seed[1970],seed[2979],seed[1357],seed[3644],seed[69],seed[4019],seed[2868],seed[1032],seed[577],seed[2203],seed[3658],seed[3568],seed[2389],seed[798],seed[417],seed[1333],seed[2068],seed[349],seed[1210],seed[489],seed[541],seed[2506],seed[971],seed[2408],seed[3602],seed[3524],seed[3196],seed[4049],seed[1875],seed[1253],seed[2667],seed[253],seed[1633],seed[302],seed[658],seed[681],seed[2308],seed[1764],seed[2637],seed[2351],seed[4060],seed[1377],seed[2027],seed[1298],seed[3688],seed[1903],seed[877],seed[2918],seed[3883],seed[2668],seed[436],seed[1587],seed[2982],seed[8],seed[2686],seed[3104],seed[2991],seed[2272],seed[3183],seed[2011],seed[365],seed[2999],seed[2948],seed[3572],seed[2165],seed[3533],seed[101],seed[1675],seed[1818],seed[814],seed[2321],seed[2022],seed[1219],seed[1543],seed[1236],seed[2398],seed[691],seed[1250],seed[839],seed[2664],seed[328],seed[1827],seed[313],seed[2429],seed[476],seed[1206],seed[2066],seed[230],seed[2117],seed[2857],seed[2849],seed[308],seed[534],seed[3784],seed[3432],seed[3212],seed[2493],seed[2467],seed[516],seed[3731],seed[578],seed[4021],seed[704],seed[460],seed[4034],seed[2738],seed[3258],seed[486],seed[752],seed[4082],seed[1862],seed[3456],seed[3168],seed[2768],seed[729],seed[2020],seed[3162],seed[3749],seed[2990],seed[1872],seed[1865],seed[376],seed[3384],seed[1503],seed[51],seed[2050],seed[1235],seed[425],seed[2485],seed[1386],seed[3845],seed[723],seed[1419],seed[804],seed[925],seed[1292],seed[2908],seed[3106],seed[256],seed[3564],seed[3917],seed[3092],seed[1525],seed[3994],seed[1312],seed[1402],seed[1802],seed[1489],seed[1696],seed[791],seed[3484],seed[199],seed[2995],seed[523],seed[3203],seed[2961],seed[220],seed[369],seed[3844],seed[2603],seed[165],seed[3216],seed[1759],seed[2093],seed[968],seed[215],seed[2481],seed[3531],seed[1632],seed[2984],seed[869],seed[2943],seed[3872],seed[2301],seed[12],seed[3767],seed[1958],seed[2670],seed[2771],seed[3346],seed[3640],seed[440],seed[3504],seed[186],seed[973],seed[2082],seed[3507],seed[1147],seed[1588],seed[2430],seed[935],seed[1189],seed[571],seed[1710],seed[3370],seed[743],seed[3809],seed[524],seed[397],seed[2407],seed[408],seed[1749],seed[2595],seed[595],seed[2314],seed[3772],seed[4093],seed[1405],seed[1897],seed[4006],seed[2568],seed[1829],seed[3894],seed[2919],seed[3285],seed[1432],seed[818],seed[2907],seed[404],seed[2711],seed[3026],seed[1861],seed[2310],seed[279],seed[3436],seed[1231],seed[211],seed[950],seed[1168],seed[332],seed[3340],seed[3388],seed[3171],seed[875],seed[1001],seed[3881],seed[1957],seed[1655],seed[42],seed[1420],seed[3007],seed[954],seed[49],seed[1596],seed[1777],seed[2873],seed[1309],seed[1146],seed[1262],seed[2780],seed[1499],seed[2897],seed[3093],seed[1563],seed[692],seed[3552],seed[2789],seed[2284],seed[166],seed[932],seed[2001],seed[2441],seed[424],seed[1247],seed[507],seed[1527],seed[1317],seed[1845],seed[3402],seed[2813],seed[2249],seed[2235],seed[3976],seed[3645],seed[1797],seed[640],seed[2935],seed[2725],seed[871],seed[3647],seed[471],seed[2553],seed[188],seed[949],seed[1974],seed[1042],seed[1211],seed[1476],seed[2562],seed[1006],seed[3099],seed[2],seed[1980],seed[1014],seed[842],seed[858],seed[560],seed[92],seed[2024],seed[2197],seed[1807],seed[2268],seed[1276],seed[1992],seed[3795],seed[556],seed[1892],seed[3462],seed[1339],seed[219],seed[2424],seed[2064],seed[114],seed[2610],seed[2227],seed[2954],seed[900],seed[1786],seed[1869],seed[2376],seed[2521],seed[19],seed[1245],seed[1224],seed[824],seed[39],seed[1997],seed[226],seed[1811],seed[1203],seed[2944],seed[1506],seed[1918],seed[2132],seed[1501],seed[2374],seed[152],seed[678],seed[3841],seed[3780],seed[3024],seed[1721],seed[1659],seed[241],seed[1776],seed[3627],seed[584],seed[2947],seed[3147],seed[3904],seed[3838],seed[1431],seed[1368],seed[1238],seed[61],seed[2869],seed[784],seed[553],seed[1899],seed[2448],seed[2015],seed[2060],seed[1084],seed[2054],seed[1604],seed[2455],seed[2309],seed[1681],seed[2150],seed[3989],seed[3320],seed[748],seed[1719],seed[1589],seed[992],seed[2953],seed[526],seed[3363],seed[3473],seed[3797],seed[1606],seed[2341],seed[4023],seed[3266],seed[3464],seed[3001],seed[3016],seed[667],seed[3313],seed[481],seed[633],seed[461],seed[4085],seed[2814],seed[1682],seed[20],seed[1272],seed[4092],seed[3996],seed[1474],seed[3421],seed[682],seed[1303],seed[3839],seed[3069],seed[537],seed[3479],seed[3133],seed[1096],seed[1263],seed[3136],seed[786],seed[3908],seed[549],seed[2864],seed[945],seed[768],seed[1566],seed[4011],seed[1856],seed[2684],seed[2119],seed[3262],seed[3933],seed[88],seed[893],seed[3758],seed[2618],seed[3332],seed[3103],seed[3950],seed[3405],seed[2271],seed[603],seed[3469],seed[2639],seed[1541],seed[2625],seed[344],seed[208],seed[3115],seed[3505],seed[2075],seed[1852],seed[379],seed[3859],seed[1578],seed[705],seed[1442],seed[2223],seed[304],seed[990],seed[1951],seed[1182],seed[2884],seed[3803],seed[143],seed[2665],seed[2804],seed[2547],seed[1979],seed[1025],seed[295],seed[2940],seed[840],seed[24],seed[1417],seed[1985],seed[3051],seed[141],seed[4008],seed[1195],seed[46],seed[1311],seed[1024],seed[1322],seed[969],seed[29],seed[2089],seed[2576],seed[2386],seed[698],seed[299],seed[754],seed[835],seed[1733],seed[112],seed[2957],seed[111],seed[323],seed[1271],seed[3261],seed[3497],seed[2342],seed[3800],seed[1495],seed[3004],seed[1075],seed[70],seed[1082],seed[117],seed[1409],seed[674],seed[3003],seed[2764],seed[2525],seed[2805],seed[2735],seed[1260],seed[3097],seed[663],seed[2199],seed[2034],seed[3459],seed[1593],seed[2882],seed[451],seed[4028],seed[802],seed[2355],seed[3457],seed[479],seed[3170],seed[706],seed[1049],seed[562],seed[757],seed[811],seed[3264],seed[1374],seed[2890],seed[1947],seed[2047],seed[3467],seed[392],seed[3761],seed[1074],seed[583],seed[1652],seed[1619],seed[2077],seed[2927],seed[3139],seed[445],seed[3977],seed[2709],seed[2803],seed[653],seed[1779],seed[2273],seed[1121],seed[175],seed[3922],seed[1510],seed[3164],seed[3736],seed[3478],seed[4065],seed[3199],seed[2615],seed[3751],seed[243],seed[4061],seed[3936],seed[1241],seed[2283],seed[619],seed[2878],seed[58],seed[1498],seed[4062],seed[1226],seed[776],seed[3878],seed[963],seed[183],seed[2096],seed[3601],seed[3327],seed[1403],seed[419],seed[733],seed[3454],seed[2827],seed[1022],seed[1880],seed[4048],seed[3991],seed[1799],seed[2841],seed[2599],seed[3987],seed[1440],seed[2695],seed[1343],seed[2536],seed[2538],seed[3906],seed[3903],seed[599],seed[2147],seed[2928],seed[3237],seed[518],seed[2008],seed[3124],seed[1701],seed[2167],seed[3949],seed[2682],seed[4058],seed[3889],seed[2035],seed[1393],seed[1728],seed[3810],seed[697],seed[3792],seed[805],seed[880],seed[2516],seed[545],seed[3389],seed[3570],seed[1978],seed[744],seed[1065],seed[1003],seed[2345],seed[1416],seed[3041],seed[659],seed[3033],seed[1021],seed[1870],seed[3480],seed[724],seed[521],seed[2874],seed[31],seed[1111],seed[564],seed[890],seed[825],seed[1944],seed[2777],seed[2741],seed[987],seed[657],seed[1427],seed[261],seed[639],seed[3495],seed[483],seed[3545],seed[116],seed[3774],seed[103],seed[3567],seed[2102],seed[1663],seed[3166],seed[3485],seed[3135],seed[3958],seed[3060],seed[2699],seed[2236],seed[2659],seed[1165],seed[148],seed[747],seed[434],seed[326],seed[2081],seed[3367],seed[3635],seed[1855],seed[1052],seed[856],seed[2337],seed[1522],seed[2619],seed[2146],seed[2561],seed[1557],seed[2023],seed[3716],seed[3945],seed[868],seed[2131],seed[1002],seed[3127],seed[1394],seed[2021],seed[3014],seed[1509],seed[3571],seed[2951],seed[2416],seed[2100],seed[2518],seed[2330],seed[2266],seed[896],seed[3948],seed[4027],seed[469],seed[1274],seed[3951],seed[1736],seed[2934],seed[277],seed[2955],seed[1819],seed[3895],seed[3373],seed[3494],seed[2009],seed[3689],seed[1467],seed[2895],seed[2248],seed[28],seed[1591],seed[1044],seed[210],seed[200],seed[1130],seed[3931],seed[1621],seed[2924],seed[1766],seed[509],seed[318],seed[1611],seed[4000],seed[1178],seed[3002],seed[3823],seed[3008],seed[3091],seed[1998],seed[1584],seed[1585],seed[2405],seed[1464],seed[632],seed[3870],seed[3757],seed[517],seed[2532],seed[1914],seed[2434],seed[1293],seed[1360],seed[1005],seed[478],seed[3760],seed[350],seed[1553],seed[1887],seed[449],seed[1194],seed[1669],seed[1067],seed[1056],seed[3413],seed[2906],seed[2811],seed[3152],seed[1039],seed[2612],seed[273],seed[2014],seed[2893],seed[922],seed[894],seed[1295],seed[3201],seed[44],seed[3597],seed[2721],seed[530],seed[2224],seed[446],seed[1127],seed[590],seed[1347],seed[316],seed[1204],seed[3530],seed[3998],seed[2140],seed[1208],seed[1592],seed[3177],seed[1949],seed[3491],seed[3296],seed[2238],seed[3218],seed[1847],seed[3848],seed[3294],seed[3409],seed[3461],seed[2976],seed[3188],seed[1688],seed[2524],seed[1012],seed[2316],seed[212],seed[938],seed[3291],seed[162],seed[3474],seed[1905],seed[3930],seed[1693],seed[122],seed[2860],seed[18],seed[1674],seed[3431],seed[353],seed[2329],seed[1485],seed[1603],seed[82],seed[1329],seed[3700],seed[1991],seed[1191],seed[1062],seed[2458],seed[2130],seed[2335],seed[3891],seed[21],seed[1546],seed[1536],seed[3347],seed[96],seed[3125],seed[2844],seed[2306],seed[2791],seed[3141],seed[687],seed[1400],seed[3455],seed[4005],seed[4001],seed[3603],seed[1441],seed[1954],seed[1275],seed[3956],seed[1645],seed[3017],seed[3290],seed[1144],seed[2902],seed[3312],seed[1977],seed[3223],seed[225],seed[2802],seed[3911],seed[2700],seed[569],seed[3306],seed[2029],seed[3849],seed[1877],seed[4044],seed[242],seed[3543],seed[3615],seed[498],seed[3526],seed[1043],seed[3050],seed[3867],seed[2913],seed[468],seed[1214],seed[2317],seed[2715],seed[936],seed[2152],seed[259],seed[3509],seed[2563],seed[3733],seed[1981],seed[1995],seed[3292],seed[3899],seed[3078],seed[2438],seed[3663],seed[1791],seed[1834],seed[1456],seed[303],seed[2067],seed[1907],seed[2819],seed[327],seed[1735],seed[3475],seed[1643],seed[2118],seed[2828],seed[3273],seed[3831],seed[2540],seed[146],seed[712],seed[1488],seed[1041],seed[669],seed[236],seed[248],seed[4004],seed[472],seed[3065],seed[385],seed[3591],seed[3159],seed[63],seed[966],seed[10],seed[3422],seed[2149],seed[3734],seed[3349],seed[3038],seed[2231],seed[1324],seed[2210],seed[2362],seed[1982],seed[2751],seed[565],seed[1487],seed[666],seed[2797],seed[2905],seed[3156],seed[2333],seed[1323],seed[180],seed[891],seed[1972],seed[3149],seed[100],seed[770],seed[2262],seed[1894],seed[2477],seed[515],seed[3310],seed[1837],seed[1821],seed[1756],seed[2511],seed[3837],seed[1774],seed[1874],seed[3999],seed[1504],seed[1934],seed[1222],seed[3244],seed[1812],seed[4075],seed[3245],seed[1114],seed[1975],seed[2270],seed[3446],seed[2694],seed[1966],seed[194],seed[1822],seed[2909],seed[158],seed[23],seed[2463],seed[3985],seed[3593],seed[1484],seed[221],seed[1909],seed[3589],seed[3990],seed[2259],seed[552],seed[2137],seed[2417],seed[139],seed[1858],seed[30],seed[3379],seed[3909],seed[3353],seed[3661],seed[919],seed[314],seed[3255],seed[93],seed[94],seed[2263],seed[2439],seed[3225],seed[1363],seed[3783],seed[458],seed[2762],seed[1131],seed[1389],seed[2313],seed[310],seed[1851],seed[3637],seed[3126],seed[2628],seed[2155],seed[3808],seed[37],seed[3673],seed[3633],seed[3054],seed[2418],seed[841],seed[3668],seed[1355],seed[1515],seed[3039],seed[1714],seed[3960],seed[2593],seed[912],seed[1330],seed[3085],seed[1428],seed[409],seed[403],seed[915],seed[1267],seed[1904],seed[2824],seed[1050],seed[3655],seed[1784],seed[671],seed[2688],seed[3653],seed[3350],seed[3020],seed[2304],seed[844],seed[466],seed[3271],seed[206],seed[1846],seed[1077],seed[3935],seed[3779],seed[216],seed[40],seed[753],seed[622],seed[2190],seed[2332],seed[495],seed[1613],seed[735],seed[2208],seed[2774],seed[513],seed[1457],seed[3755],seed[977],seed[3123],seed[3538],seed[2614],seed[1900],seed[1703],seed[3967],seed[1451],seed[1265],seed[3798],seed[3660],seed[1029],seed[2710],seed[1149],seed[90],seed[2298],seed[3687],seed[3437],seed[2978],seed[2733],seed[1744],seed[3034],seed[280],seed[1864],seed[1512],seed[547],seed[3821],seed[99],seed[429],seed[2276],seed[1524],seed[1233],seed[1910],seed[3836],seed[3321],seed[1685],seed[1358],seed[3665],seed[1229],seed[3143],seed[2300],seed[3068],seed[1550],seed[1554],seed[2973],seed[3675],seed[2013],seed[1156],seed[2977],seed[2649],seed[1070],seed[3807],seed[2127],seed[284],seed[2475],seed[2696],seed[1508],seed[1469],seed[3438],seed[879],seed[2039],seed[366],seed[3723],seed[3997],seed[1540],seed[2136],seed[3406],seed[1388],seed[2491],seed[718],seed[3852],seed[1346],seed[3793],seed[831],seed[3331],seed[4002],seed[2838],seed[1083],seed[1939],seed[266],seed[3280],seed[106],seed[2312],seed[921],seed[2914],seed[956],seed[2296],seed[1255],seed[1867],seed[159],seed[937],seed[1545],seed[1810],seed[2187],seed[3448],seed[3885],seed[2207],seed[3879],seed[3847],seed[3943],seed[2324],seed[156],seed[1935],seed[2885],seed[3163],seed[2656],seed[2053],seed[2754],seed[854],seed[2396],seed[3443],seed[1391],seed[700],seed[3840],seed[1300],seed[853],seed[2171],seed[1422],seed[3611],seed[567],seed[2279],seed[1151],seed[1397],seed[3299],seed[2969],seed[1101],seed[907],seed[1369],seed[3302],seed[3801],seed[4080],seed[2815],seed[245],seed[1994],seed[2178],seed[2290],seed[3305],seed[1636],seed[1406],seed[2833],seed[2206],seed[1729],seed[4022],seed[2120],seed[3073],seed[2359],seed[866],seed[872],seed[2242],seed[684],seed[2745],seed[2703],seed[2956],seed[336],seed[1152],seed[3359],seed[2225],seed[2717],seed[766],seed[2452],seed[3995],seed[2151],seed[625],seed[3714],seed[1028],seed[3510],seed[278],seed[337],seed[3101],seed[4051],seed[1354],seed[2125],seed[431],seed[1412],seed[1787],seed[1199],seed[3874],seed[902],seed[2031],seed[2706],seed[1739],seed[2636],seed[2830],seed[2915],seed[3866],seed[2886],seed[721],seed[3659],seed[1294],seed[2468],seed[60],seed[1941],seed[235],seed[1244],seed[430],seed[2320],seed[2911],seed[319],seed[2965],seed[1332],seed[1668],seed[427],seed[1745],seed[2443],seed[604],seed[3129],seed[131],seed[2846],seed[2461],seed[1249],seed[2671],seed[1026],seed[258],seed[926],seed[1754],seed[3098],seed[1450],seed[50],seed[3449],seed[470],seed[1308],seed[2580],seed[1390],seed[170],seed[2597],seed[3692],seed[2801],seed[1727],seed[2613],seed[1023],seed[3062],seed[548],seed[2980],seed[351],seed[3566],seed[2212],seed[1110],seed[3090],seed[3501],seed[2749],seed[2447],seed[3499],seed[538],seed[2596],seed[2221],seed[808],seed[1608],seed[315],seed[3391],seed[3514],seed[2507],seed[2623],seed[3077],seed[3374],seed[1171],seed[1930],seed[4074],seed[1107],seed[2528],seed[3992],seed[3214],seed[393],seed[675],seed[3013],seed[594],seed[1018],seed[3833],seed[3677],seed[694],seed[1282],seed[1559],seed[2912],seed[3898],seed[4081],seed[2142],seed[2926],seed[693]}),
        .cross_prob(cross_prob),
        .codeword(codeword16),
        .received(received16)
        );
    
//    bsc bsc1(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed1),
//        .cross_prob(cross_prob),
//        .codeword(codeword1),
//        .received(received1)
//        );
    
//    bsc bsc2(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed2),
//        .cross_prob(cross_prob),
//        .codeword(codeword2),
//        .received(received2)
//        );
        
//    bsc bsc3(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed3),
//        .cross_prob(cross_prob),
//        .codeword(codeword3),
//        .received(received3)
//        );
    
//    bsc bsc4(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed4),
//        .cross_prob(cross_prob),
//        .codeword(codeword4),
//        .received(received4)
//        );
    
//    bsc bsc5(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed5),
//        .cross_prob(cross_prob),
//        .codeword(codeword5),
//        .received(received5)
//        );
    
//    bsc bsc6(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed6),
//        .cross_prob(cross_prob),
//        .codeword(codeword6),
//        .received(received6)
//        );
    
//    bsc bsc7(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed7),
//        .cross_prob(cross_prob),
//        .codeword(codeword7),
//        .received(received7)
//        );
        
//    bsc bsc8(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed8),
//        .cross_prob(cross_prob),
//        .codeword(codeword8),
//        .received(received8)
//        );
    
//    bsc bsc9(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed9),
//        .cross_prob(cross_prob),
//        .codeword(codeword9),
//        .received(received9)
//        );
    
//    bsc bsc10(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed10),
//        .cross_prob(cross_prob),
//        .codeword(codeword10),
//        .received(received10)
//        );
    
//    bsc bsc11(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed11),
//        .cross_prob(cross_prob),
//        .codeword(codeword11),
//        .received(received11)
//        );
    
//    bsc bsc12(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed12),
//        .cross_prob(cross_prob),
//        .codeword(codeword12),
//        .received(received12)
//        );
    
//    bsc bsc13(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed13),
//        .cross_prob(cross_prob),
//        .codeword(codeword13),
//        .received(received13)
//        );
    
//    bsc bsc14(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed14),
//        .cross_prob(cross_prob),
//        .codeword(codeword14),
//        .received(received14)
//        );
    
//    bsc bsc15(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed15),
//        .cross_prob(cross_prob),
//        .codeword(codeword15),
//        .received(received15)
//        );
    
//    bsc bsc16(
//        .clk(clk),
//        .reset(reset),
//        .seed(seed16),
//        .cross_prob(cross_prob),
//        .codeword(codeword16),
//        .received(received16)
//        );
    
    
endmodule